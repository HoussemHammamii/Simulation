`timescale 1 ns/1 ps

module MeshOfTree(
     clock
   , conf
   , reset
   , address
   , data
   , inpads_top
   , inpads_right
   , inpads_bottom
   , inpads_left
   , outpads_top
   , outpads_right
   , outpads_bottom
   , outpads_left
  );


input   clock;
wire clock;
input   conf;
wire conf;
input   reset;
wire reset;
input   [14:0] address;
wire [14:0] address;
input   [7:0] data;
wire [7:0] data;
input   [7:0] inpads_top;
wire [7:0] inpads_top;
input   [7:0] inpads_right;
wire [7:0] inpads_right;
input   [7:0] inpads_bottom;
wire [7:0] inpads_bottom;
input   [7:0] inpads_left;
wire [7:0] inpads_left;
output  [7:0] outpads_top;
wire [7:0] outpads_top;
output  [7:0] outpads_right;
wire [7:0] outpads_right;
output  [7:0] outpads_bottom;
wire [7:0] outpads_bottom;
output  [7:0] outpads_left;
wire [7:0] outpads_left;

wire wire_in_cluster_sb_BL_0_0;
wire wire_in_cluster_sb_BL_0_1;
wire wire_in_cluster_sb_BL_0_10;
wire wire_in_cluster_sb_BL_0_11;
wire wire_in_cluster_sb_BL_0_12;
wire wire_in_cluster_sb_BL_0_13;
wire wire_in_cluster_sb_BL_0_14;
wire wire_in_cluster_sb_BL_0_15;
wire wire_in_cluster_sb_BL_0_2;
wire wire_in_cluster_sb_BL_0_3;
wire wire_in_cluster_sb_BL_0_4;
wire wire_in_cluster_sb_BL_0_5;
wire wire_in_cluster_sb_BL_0_6;
wire wire_in_cluster_sb_BL_0_7;
wire wire_in_cluster_sb_BL_0_8;
wire wire_in_cluster_sb_BL_0_9;
wire wire_in_cluster_sb_BL_10_0;
wire wire_in_cluster_sb_BL_10_1;
wire wire_in_cluster_sb_BL_10_10;
wire wire_in_cluster_sb_BL_10_11;
wire wire_in_cluster_sb_BL_10_12;
wire wire_in_cluster_sb_BL_10_13;
wire wire_in_cluster_sb_BL_10_14;
wire wire_in_cluster_sb_BL_10_15;
wire wire_in_cluster_sb_BL_10_2;
wire wire_in_cluster_sb_BL_10_3;
wire wire_in_cluster_sb_BL_10_4;
wire wire_in_cluster_sb_BL_10_5;
wire wire_in_cluster_sb_BL_10_6;
wire wire_in_cluster_sb_BL_10_7;
wire wire_in_cluster_sb_BL_10_8;
wire wire_in_cluster_sb_BL_10_9;
wire wire_in_cluster_sb_BL_11_0;
wire wire_in_cluster_sb_BL_11_1;
wire wire_in_cluster_sb_BL_11_10;
wire wire_in_cluster_sb_BL_11_11;
wire wire_in_cluster_sb_BL_11_12;
wire wire_in_cluster_sb_BL_11_13;
wire wire_in_cluster_sb_BL_11_14;
wire wire_in_cluster_sb_BL_11_15;
wire wire_in_cluster_sb_BL_11_2;
wire wire_in_cluster_sb_BL_11_3;
wire wire_in_cluster_sb_BL_11_4;
wire wire_in_cluster_sb_BL_11_5;
wire wire_in_cluster_sb_BL_11_6;
wire wire_in_cluster_sb_BL_11_7;
wire wire_in_cluster_sb_BL_11_8;
wire wire_in_cluster_sb_BL_11_9;
wire wire_in_cluster_sb_BL_12_0;
wire wire_in_cluster_sb_BL_12_1;
wire wire_in_cluster_sb_BL_12_10;
wire wire_in_cluster_sb_BL_12_11;
wire wire_in_cluster_sb_BL_12_12;
wire wire_in_cluster_sb_BL_12_13;
wire wire_in_cluster_sb_BL_12_14;
wire wire_in_cluster_sb_BL_12_15;
wire wire_in_cluster_sb_BL_12_2;
wire wire_in_cluster_sb_BL_12_3;
wire wire_in_cluster_sb_BL_12_4;
wire wire_in_cluster_sb_BL_12_5;
wire wire_in_cluster_sb_BL_12_6;
wire wire_in_cluster_sb_BL_12_7;
wire wire_in_cluster_sb_BL_12_8;
wire wire_in_cluster_sb_BL_12_9;
wire wire_in_cluster_sb_BL_13_0;
wire wire_in_cluster_sb_BL_13_1;
wire wire_in_cluster_sb_BL_13_10;
wire wire_in_cluster_sb_BL_13_11;
wire wire_in_cluster_sb_BL_13_12;
wire wire_in_cluster_sb_BL_13_13;
wire wire_in_cluster_sb_BL_13_14;
wire wire_in_cluster_sb_BL_13_15;
wire wire_in_cluster_sb_BL_13_2;
wire wire_in_cluster_sb_BL_13_3;
wire wire_in_cluster_sb_BL_13_4;
wire wire_in_cluster_sb_BL_13_5;
wire wire_in_cluster_sb_BL_13_6;
wire wire_in_cluster_sb_BL_13_7;
wire wire_in_cluster_sb_BL_13_8;
wire wire_in_cluster_sb_BL_13_9;
wire wire_in_cluster_sb_BL_14_0;
wire wire_in_cluster_sb_BL_14_1;
wire wire_in_cluster_sb_BL_14_10;
wire wire_in_cluster_sb_BL_14_11;
wire wire_in_cluster_sb_BL_14_12;
wire wire_in_cluster_sb_BL_14_13;
wire wire_in_cluster_sb_BL_14_14;
wire wire_in_cluster_sb_BL_14_15;
wire wire_in_cluster_sb_BL_14_2;
wire wire_in_cluster_sb_BL_14_3;
wire wire_in_cluster_sb_BL_14_4;
wire wire_in_cluster_sb_BL_14_5;
wire wire_in_cluster_sb_BL_14_6;
wire wire_in_cluster_sb_BL_14_7;
wire wire_in_cluster_sb_BL_14_8;
wire wire_in_cluster_sb_BL_14_9;
wire wire_in_cluster_sb_BL_15_0;
wire wire_in_cluster_sb_BL_15_1;
wire wire_in_cluster_sb_BL_15_10;
wire wire_in_cluster_sb_BL_15_11;
wire wire_in_cluster_sb_BL_15_12;
wire wire_in_cluster_sb_BL_15_13;
wire wire_in_cluster_sb_BL_15_14;
wire wire_in_cluster_sb_BL_15_15;
wire wire_in_cluster_sb_BL_15_2;
wire wire_in_cluster_sb_BL_15_3;
wire wire_in_cluster_sb_BL_15_4;
wire wire_in_cluster_sb_BL_15_5;
wire wire_in_cluster_sb_BL_15_6;
wire wire_in_cluster_sb_BL_15_7;
wire wire_in_cluster_sb_BL_15_8;
wire wire_in_cluster_sb_BL_15_9;
wire wire_in_cluster_sb_BL_1_0;
wire wire_in_cluster_sb_BL_1_1;
wire wire_in_cluster_sb_BL_1_10;
wire wire_in_cluster_sb_BL_1_11;
wire wire_in_cluster_sb_BL_1_12;
wire wire_in_cluster_sb_BL_1_13;
wire wire_in_cluster_sb_BL_1_14;
wire wire_in_cluster_sb_BL_1_15;
wire wire_in_cluster_sb_BL_1_2;
wire wire_in_cluster_sb_BL_1_3;
wire wire_in_cluster_sb_BL_1_4;
wire wire_in_cluster_sb_BL_1_5;
wire wire_in_cluster_sb_BL_1_6;
wire wire_in_cluster_sb_BL_1_7;
wire wire_in_cluster_sb_BL_1_8;
wire wire_in_cluster_sb_BL_1_9;
wire wire_in_cluster_sb_BL_2_0;
wire wire_in_cluster_sb_BL_2_1;
wire wire_in_cluster_sb_BL_2_10;
wire wire_in_cluster_sb_BL_2_11;
wire wire_in_cluster_sb_BL_2_12;
wire wire_in_cluster_sb_BL_2_13;
wire wire_in_cluster_sb_BL_2_14;
wire wire_in_cluster_sb_BL_2_15;
wire wire_in_cluster_sb_BL_2_2;
wire wire_in_cluster_sb_BL_2_3;
wire wire_in_cluster_sb_BL_2_4;
wire wire_in_cluster_sb_BL_2_5;
wire wire_in_cluster_sb_BL_2_6;
wire wire_in_cluster_sb_BL_2_7;
wire wire_in_cluster_sb_BL_2_8;
wire wire_in_cluster_sb_BL_2_9;
wire wire_in_cluster_sb_BL_3_0;
wire wire_in_cluster_sb_BL_3_1;
wire wire_in_cluster_sb_BL_3_10;
wire wire_in_cluster_sb_BL_3_11;
wire wire_in_cluster_sb_BL_3_12;
wire wire_in_cluster_sb_BL_3_13;
wire wire_in_cluster_sb_BL_3_14;
wire wire_in_cluster_sb_BL_3_15;
wire wire_in_cluster_sb_BL_3_2;
wire wire_in_cluster_sb_BL_3_3;
wire wire_in_cluster_sb_BL_3_4;
wire wire_in_cluster_sb_BL_3_5;
wire wire_in_cluster_sb_BL_3_6;
wire wire_in_cluster_sb_BL_3_7;
wire wire_in_cluster_sb_BL_3_8;
wire wire_in_cluster_sb_BL_3_9;
wire wire_in_cluster_sb_BL_4_0;
wire wire_in_cluster_sb_BL_4_1;
wire wire_in_cluster_sb_BL_4_10;
wire wire_in_cluster_sb_BL_4_11;
wire wire_in_cluster_sb_BL_4_12;
wire wire_in_cluster_sb_BL_4_13;
wire wire_in_cluster_sb_BL_4_14;
wire wire_in_cluster_sb_BL_4_15;
wire wire_in_cluster_sb_BL_4_2;
wire wire_in_cluster_sb_BL_4_3;
wire wire_in_cluster_sb_BL_4_4;
wire wire_in_cluster_sb_BL_4_5;
wire wire_in_cluster_sb_BL_4_6;
wire wire_in_cluster_sb_BL_4_7;
wire wire_in_cluster_sb_BL_4_8;
wire wire_in_cluster_sb_BL_4_9;
wire wire_in_cluster_sb_BL_5_0;
wire wire_in_cluster_sb_BL_5_1;
wire wire_in_cluster_sb_BL_5_10;
wire wire_in_cluster_sb_BL_5_11;
wire wire_in_cluster_sb_BL_5_12;
wire wire_in_cluster_sb_BL_5_13;
wire wire_in_cluster_sb_BL_5_14;
wire wire_in_cluster_sb_BL_5_15;
wire wire_in_cluster_sb_BL_5_2;
wire wire_in_cluster_sb_BL_5_3;
wire wire_in_cluster_sb_BL_5_4;
wire wire_in_cluster_sb_BL_5_5;
wire wire_in_cluster_sb_BL_5_6;
wire wire_in_cluster_sb_BL_5_7;
wire wire_in_cluster_sb_BL_5_8;
wire wire_in_cluster_sb_BL_5_9;
wire wire_in_cluster_sb_BL_6_0;
wire wire_in_cluster_sb_BL_6_1;
wire wire_in_cluster_sb_BL_6_10;
wire wire_in_cluster_sb_BL_6_11;
wire wire_in_cluster_sb_BL_6_12;
wire wire_in_cluster_sb_BL_6_13;
wire wire_in_cluster_sb_BL_6_14;
wire wire_in_cluster_sb_BL_6_15;
wire wire_in_cluster_sb_BL_6_2;
wire wire_in_cluster_sb_BL_6_3;
wire wire_in_cluster_sb_BL_6_4;
wire wire_in_cluster_sb_BL_6_5;
wire wire_in_cluster_sb_BL_6_6;
wire wire_in_cluster_sb_BL_6_7;
wire wire_in_cluster_sb_BL_6_8;
wire wire_in_cluster_sb_BL_6_9;
wire wire_in_cluster_sb_BL_7_0;
wire wire_in_cluster_sb_BL_7_1;
wire wire_in_cluster_sb_BL_7_10;
wire wire_in_cluster_sb_BL_7_11;
wire wire_in_cluster_sb_BL_7_12;
wire wire_in_cluster_sb_BL_7_13;
wire wire_in_cluster_sb_BL_7_14;
wire wire_in_cluster_sb_BL_7_15;
wire wire_in_cluster_sb_BL_7_2;
wire wire_in_cluster_sb_BL_7_3;
wire wire_in_cluster_sb_BL_7_4;
wire wire_in_cluster_sb_BL_7_5;
wire wire_in_cluster_sb_BL_7_6;
wire wire_in_cluster_sb_BL_7_7;
wire wire_in_cluster_sb_BL_7_8;
wire wire_in_cluster_sb_BL_7_9;
wire wire_in_cluster_sb_BL_8_0;
wire wire_in_cluster_sb_BL_8_1;
wire wire_in_cluster_sb_BL_8_10;
wire wire_in_cluster_sb_BL_8_11;
wire wire_in_cluster_sb_BL_8_12;
wire wire_in_cluster_sb_BL_8_13;
wire wire_in_cluster_sb_BL_8_14;
wire wire_in_cluster_sb_BL_8_15;
wire wire_in_cluster_sb_BL_8_2;
wire wire_in_cluster_sb_BL_8_3;
wire wire_in_cluster_sb_BL_8_4;
wire wire_in_cluster_sb_BL_8_5;
wire wire_in_cluster_sb_BL_8_6;
wire wire_in_cluster_sb_BL_8_7;
wire wire_in_cluster_sb_BL_8_8;
wire wire_in_cluster_sb_BL_8_9;
wire wire_in_cluster_sb_BL_9_0;
wire wire_in_cluster_sb_BL_9_1;
wire wire_in_cluster_sb_BL_9_10;
wire wire_in_cluster_sb_BL_9_11;
wire wire_in_cluster_sb_BL_9_12;
wire wire_in_cluster_sb_BL_9_13;
wire wire_in_cluster_sb_BL_9_14;
wire wire_in_cluster_sb_BL_9_15;
wire wire_in_cluster_sb_BL_9_2;
wire wire_in_cluster_sb_BL_9_3;
wire wire_in_cluster_sb_BL_9_4;
wire wire_in_cluster_sb_BL_9_5;
wire wire_in_cluster_sb_BL_9_6;
wire wire_in_cluster_sb_BL_9_7;
wire wire_in_cluster_sb_BL_9_8;
wire wire_in_cluster_sb_BL_9_9;
wire wire_in_cluster_sb_BR_0_0;
wire wire_in_cluster_sb_BR_0_1;
wire wire_in_cluster_sb_BR_0_10;
wire wire_in_cluster_sb_BR_0_11;
wire wire_in_cluster_sb_BR_0_12;
wire wire_in_cluster_sb_BR_0_13;
wire wire_in_cluster_sb_BR_0_14;
wire wire_in_cluster_sb_BR_0_15;
wire wire_in_cluster_sb_BR_0_2;
wire wire_in_cluster_sb_BR_0_3;
wire wire_in_cluster_sb_BR_0_4;
wire wire_in_cluster_sb_BR_0_5;
wire wire_in_cluster_sb_BR_0_6;
wire wire_in_cluster_sb_BR_0_7;
wire wire_in_cluster_sb_BR_0_8;
wire wire_in_cluster_sb_BR_0_9;
wire wire_in_cluster_sb_BR_10_0;
wire wire_in_cluster_sb_BR_10_1;
wire wire_in_cluster_sb_BR_10_10;
wire wire_in_cluster_sb_BR_10_11;
wire wire_in_cluster_sb_BR_10_12;
wire wire_in_cluster_sb_BR_10_13;
wire wire_in_cluster_sb_BR_10_14;
wire wire_in_cluster_sb_BR_10_15;
wire wire_in_cluster_sb_BR_10_2;
wire wire_in_cluster_sb_BR_10_3;
wire wire_in_cluster_sb_BR_10_4;
wire wire_in_cluster_sb_BR_10_5;
wire wire_in_cluster_sb_BR_10_6;
wire wire_in_cluster_sb_BR_10_7;
wire wire_in_cluster_sb_BR_10_8;
wire wire_in_cluster_sb_BR_10_9;
wire wire_in_cluster_sb_BR_11_0;
wire wire_in_cluster_sb_BR_11_1;
wire wire_in_cluster_sb_BR_11_10;
wire wire_in_cluster_sb_BR_11_11;
wire wire_in_cluster_sb_BR_11_12;
wire wire_in_cluster_sb_BR_11_13;
wire wire_in_cluster_sb_BR_11_14;
wire wire_in_cluster_sb_BR_11_15;
wire wire_in_cluster_sb_BR_11_2;
wire wire_in_cluster_sb_BR_11_3;
wire wire_in_cluster_sb_BR_11_4;
wire wire_in_cluster_sb_BR_11_5;
wire wire_in_cluster_sb_BR_11_6;
wire wire_in_cluster_sb_BR_11_7;
wire wire_in_cluster_sb_BR_11_8;
wire wire_in_cluster_sb_BR_11_9;
wire wire_in_cluster_sb_BR_12_0;
wire wire_in_cluster_sb_BR_12_1;
wire wire_in_cluster_sb_BR_12_10;
wire wire_in_cluster_sb_BR_12_11;
wire wire_in_cluster_sb_BR_12_12;
wire wire_in_cluster_sb_BR_12_13;
wire wire_in_cluster_sb_BR_12_14;
wire wire_in_cluster_sb_BR_12_15;
wire wire_in_cluster_sb_BR_12_2;
wire wire_in_cluster_sb_BR_12_3;
wire wire_in_cluster_sb_BR_12_4;
wire wire_in_cluster_sb_BR_12_5;
wire wire_in_cluster_sb_BR_12_6;
wire wire_in_cluster_sb_BR_12_7;
wire wire_in_cluster_sb_BR_12_8;
wire wire_in_cluster_sb_BR_12_9;
wire wire_in_cluster_sb_BR_13_0;
wire wire_in_cluster_sb_BR_13_1;
wire wire_in_cluster_sb_BR_13_10;
wire wire_in_cluster_sb_BR_13_11;
wire wire_in_cluster_sb_BR_13_12;
wire wire_in_cluster_sb_BR_13_13;
wire wire_in_cluster_sb_BR_13_14;
wire wire_in_cluster_sb_BR_13_15;
wire wire_in_cluster_sb_BR_13_2;
wire wire_in_cluster_sb_BR_13_3;
wire wire_in_cluster_sb_BR_13_4;
wire wire_in_cluster_sb_BR_13_5;
wire wire_in_cluster_sb_BR_13_6;
wire wire_in_cluster_sb_BR_13_7;
wire wire_in_cluster_sb_BR_13_8;
wire wire_in_cluster_sb_BR_13_9;
wire wire_in_cluster_sb_BR_14_0;
wire wire_in_cluster_sb_BR_14_1;
wire wire_in_cluster_sb_BR_14_10;
wire wire_in_cluster_sb_BR_14_11;
wire wire_in_cluster_sb_BR_14_12;
wire wire_in_cluster_sb_BR_14_13;
wire wire_in_cluster_sb_BR_14_14;
wire wire_in_cluster_sb_BR_14_15;
wire wire_in_cluster_sb_BR_14_2;
wire wire_in_cluster_sb_BR_14_3;
wire wire_in_cluster_sb_BR_14_4;
wire wire_in_cluster_sb_BR_14_5;
wire wire_in_cluster_sb_BR_14_6;
wire wire_in_cluster_sb_BR_14_7;
wire wire_in_cluster_sb_BR_14_8;
wire wire_in_cluster_sb_BR_14_9;
wire wire_in_cluster_sb_BR_15_0;
wire wire_in_cluster_sb_BR_15_1;
wire wire_in_cluster_sb_BR_15_10;
wire wire_in_cluster_sb_BR_15_11;
wire wire_in_cluster_sb_BR_15_12;
wire wire_in_cluster_sb_BR_15_13;
wire wire_in_cluster_sb_BR_15_14;
wire wire_in_cluster_sb_BR_15_15;
wire wire_in_cluster_sb_BR_15_2;
wire wire_in_cluster_sb_BR_15_3;
wire wire_in_cluster_sb_BR_15_4;
wire wire_in_cluster_sb_BR_15_5;
wire wire_in_cluster_sb_BR_15_6;
wire wire_in_cluster_sb_BR_15_7;
wire wire_in_cluster_sb_BR_15_8;
wire wire_in_cluster_sb_BR_15_9;
wire wire_in_cluster_sb_BR_1_0;
wire wire_in_cluster_sb_BR_1_1;
wire wire_in_cluster_sb_BR_1_10;
wire wire_in_cluster_sb_BR_1_11;
wire wire_in_cluster_sb_BR_1_12;
wire wire_in_cluster_sb_BR_1_13;
wire wire_in_cluster_sb_BR_1_14;
wire wire_in_cluster_sb_BR_1_15;
wire wire_in_cluster_sb_BR_1_2;
wire wire_in_cluster_sb_BR_1_3;
wire wire_in_cluster_sb_BR_1_4;
wire wire_in_cluster_sb_BR_1_5;
wire wire_in_cluster_sb_BR_1_6;
wire wire_in_cluster_sb_BR_1_7;
wire wire_in_cluster_sb_BR_1_8;
wire wire_in_cluster_sb_BR_1_9;
wire wire_in_cluster_sb_BR_2_0;
wire wire_in_cluster_sb_BR_2_1;
wire wire_in_cluster_sb_BR_2_10;
wire wire_in_cluster_sb_BR_2_11;
wire wire_in_cluster_sb_BR_2_12;
wire wire_in_cluster_sb_BR_2_13;
wire wire_in_cluster_sb_BR_2_14;
wire wire_in_cluster_sb_BR_2_15;
wire wire_in_cluster_sb_BR_2_2;
wire wire_in_cluster_sb_BR_2_3;
wire wire_in_cluster_sb_BR_2_4;
wire wire_in_cluster_sb_BR_2_5;
wire wire_in_cluster_sb_BR_2_6;
wire wire_in_cluster_sb_BR_2_7;
wire wire_in_cluster_sb_BR_2_8;
wire wire_in_cluster_sb_BR_2_9;
wire wire_in_cluster_sb_BR_3_0;
wire wire_in_cluster_sb_BR_3_1;
wire wire_in_cluster_sb_BR_3_10;
wire wire_in_cluster_sb_BR_3_11;
wire wire_in_cluster_sb_BR_3_12;
wire wire_in_cluster_sb_BR_3_13;
wire wire_in_cluster_sb_BR_3_14;
wire wire_in_cluster_sb_BR_3_15;
wire wire_in_cluster_sb_BR_3_2;
wire wire_in_cluster_sb_BR_3_3;
wire wire_in_cluster_sb_BR_3_4;
wire wire_in_cluster_sb_BR_3_5;
wire wire_in_cluster_sb_BR_3_6;
wire wire_in_cluster_sb_BR_3_7;
wire wire_in_cluster_sb_BR_3_8;
wire wire_in_cluster_sb_BR_3_9;
wire wire_in_cluster_sb_BR_4_0;
wire wire_in_cluster_sb_BR_4_1;
wire wire_in_cluster_sb_BR_4_10;
wire wire_in_cluster_sb_BR_4_11;
wire wire_in_cluster_sb_BR_4_12;
wire wire_in_cluster_sb_BR_4_13;
wire wire_in_cluster_sb_BR_4_14;
wire wire_in_cluster_sb_BR_4_15;
wire wire_in_cluster_sb_BR_4_2;
wire wire_in_cluster_sb_BR_4_3;
wire wire_in_cluster_sb_BR_4_4;
wire wire_in_cluster_sb_BR_4_5;
wire wire_in_cluster_sb_BR_4_6;
wire wire_in_cluster_sb_BR_4_7;
wire wire_in_cluster_sb_BR_4_8;
wire wire_in_cluster_sb_BR_4_9;
wire wire_in_cluster_sb_BR_5_0;
wire wire_in_cluster_sb_BR_5_1;
wire wire_in_cluster_sb_BR_5_10;
wire wire_in_cluster_sb_BR_5_11;
wire wire_in_cluster_sb_BR_5_12;
wire wire_in_cluster_sb_BR_5_13;
wire wire_in_cluster_sb_BR_5_14;
wire wire_in_cluster_sb_BR_5_15;
wire wire_in_cluster_sb_BR_5_2;
wire wire_in_cluster_sb_BR_5_3;
wire wire_in_cluster_sb_BR_5_4;
wire wire_in_cluster_sb_BR_5_5;
wire wire_in_cluster_sb_BR_5_6;
wire wire_in_cluster_sb_BR_5_7;
wire wire_in_cluster_sb_BR_5_8;
wire wire_in_cluster_sb_BR_5_9;
wire wire_in_cluster_sb_BR_6_0;
wire wire_in_cluster_sb_BR_6_1;
wire wire_in_cluster_sb_BR_6_10;
wire wire_in_cluster_sb_BR_6_11;
wire wire_in_cluster_sb_BR_6_12;
wire wire_in_cluster_sb_BR_6_13;
wire wire_in_cluster_sb_BR_6_14;
wire wire_in_cluster_sb_BR_6_15;
wire wire_in_cluster_sb_BR_6_2;
wire wire_in_cluster_sb_BR_6_3;
wire wire_in_cluster_sb_BR_6_4;
wire wire_in_cluster_sb_BR_6_5;
wire wire_in_cluster_sb_BR_6_6;
wire wire_in_cluster_sb_BR_6_7;
wire wire_in_cluster_sb_BR_6_8;
wire wire_in_cluster_sb_BR_6_9;
wire wire_in_cluster_sb_BR_7_0;
wire wire_in_cluster_sb_BR_7_1;
wire wire_in_cluster_sb_BR_7_10;
wire wire_in_cluster_sb_BR_7_11;
wire wire_in_cluster_sb_BR_7_12;
wire wire_in_cluster_sb_BR_7_13;
wire wire_in_cluster_sb_BR_7_14;
wire wire_in_cluster_sb_BR_7_15;
wire wire_in_cluster_sb_BR_7_2;
wire wire_in_cluster_sb_BR_7_3;
wire wire_in_cluster_sb_BR_7_4;
wire wire_in_cluster_sb_BR_7_5;
wire wire_in_cluster_sb_BR_7_6;
wire wire_in_cluster_sb_BR_7_7;
wire wire_in_cluster_sb_BR_7_8;
wire wire_in_cluster_sb_BR_7_9;
wire wire_in_cluster_sb_BR_8_0;
wire wire_in_cluster_sb_BR_8_1;
wire wire_in_cluster_sb_BR_8_10;
wire wire_in_cluster_sb_BR_8_11;
wire wire_in_cluster_sb_BR_8_12;
wire wire_in_cluster_sb_BR_8_13;
wire wire_in_cluster_sb_BR_8_14;
wire wire_in_cluster_sb_BR_8_15;
wire wire_in_cluster_sb_BR_8_2;
wire wire_in_cluster_sb_BR_8_3;
wire wire_in_cluster_sb_BR_8_4;
wire wire_in_cluster_sb_BR_8_5;
wire wire_in_cluster_sb_BR_8_6;
wire wire_in_cluster_sb_BR_8_7;
wire wire_in_cluster_sb_BR_8_8;
wire wire_in_cluster_sb_BR_8_9;
wire wire_in_cluster_sb_BR_9_0;
wire wire_in_cluster_sb_BR_9_1;
wire wire_in_cluster_sb_BR_9_10;
wire wire_in_cluster_sb_BR_9_11;
wire wire_in_cluster_sb_BR_9_12;
wire wire_in_cluster_sb_BR_9_13;
wire wire_in_cluster_sb_BR_9_14;
wire wire_in_cluster_sb_BR_9_15;
wire wire_in_cluster_sb_BR_9_2;
wire wire_in_cluster_sb_BR_9_3;
wire wire_in_cluster_sb_BR_9_4;
wire wire_in_cluster_sb_BR_9_5;
wire wire_in_cluster_sb_BR_9_6;
wire wire_in_cluster_sb_BR_9_7;
wire wire_in_cluster_sb_BR_9_8;
wire wire_in_cluster_sb_BR_9_9;
wire wire_in_cluster_sb_TL_0_0;
wire wire_in_cluster_sb_TL_0_1;
wire wire_in_cluster_sb_TL_0_10;
wire wire_in_cluster_sb_TL_0_11;
wire wire_in_cluster_sb_TL_0_12;
wire wire_in_cluster_sb_TL_0_13;
wire wire_in_cluster_sb_TL_0_14;
wire wire_in_cluster_sb_TL_0_15;
wire wire_in_cluster_sb_TL_0_2;
wire wire_in_cluster_sb_TL_0_3;
wire wire_in_cluster_sb_TL_0_4;
wire wire_in_cluster_sb_TL_0_5;
wire wire_in_cluster_sb_TL_0_6;
wire wire_in_cluster_sb_TL_0_7;
wire wire_in_cluster_sb_TL_0_8;
wire wire_in_cluster_sb_TL_0_9;
wire wire_in_cluster_sb_TL_10_0;
wire wire_in_cluster_sb_TL_10_1;
wire wire_in_cluster_sb_TL_10_10;
wire wire_in_cluster_sb_TL_10_11;
wire wire_in_cluster_sb_TL_10_12;
wire wire_in_cluster_sb_TL_10_13;
wire wire_in_cluster_sb_TL_10_14;
wire wire_in_cluster_sb_TL_10_15;
wire wire_in_cluster_sb_TL_10_2;
wire wire_in_cluster_sb_TL_10_3;
wire wire_in_cluster_sb_TL_10_4;
wire wire_in_cluster_sb_TL_10_5;
wire wire_in_cluster_sb_TL_10_6;
wire wire_in_cluster_sb_TL_10_7;
wire wire_in_cluster_sb_TL_10_8;
wire wire_in_cluster_sb_TL_10_9;
wire wire_in_cluster_sb_TL_11_0;
wire wire_in_cluster_sb_TL_11_1;
wire wire_in_cluster_sb_TL_11_10;
wire wire_in_cluster_sb_TL_11_11;
wire wire_in_cluster_sb_TL_11_12;
wire wire_in_cluster_sb_TL_11_13;
wire wire_in_cluster_sb_TL_11_14;
wire wire_in_cluster_sb_TL_11_15;
wire wire_in_cluster_sb_TL_11_2;
wire wire_in_cluster_sb_TL_11_3;
wire wire_in_cluster_sb_TL_11_4;
wire wire_in_cluster_sb_TL_11_5;
wire wire_in_cluster_sb_TL_11_6;
wire wire_in_cluster_sb_TL_11_7;
wire wire_in_cluster_sb_TL_11_8;
wire wire_in_cluster_sb_TL_11_9;
wire wire_in_cluster_sb_TL_12_0;
wire wire_in_cluster_sb_TL_12_1;
wire wire_in_cluster_sb_TL_12_10;
wire wire_in_cluster_sb_TL_12_11;
wire wire_in_cluster_sb_TL_12_12;
wire wire_in_cluster_sb_TL_12_13;
wire wire_in_cluster_sb_TL_12_14;
wire wire_in_cluster_sb_TL_12_15;
wire wire_in_cluster_sb_TL_12_2;
wire wire_in_cluster_sb_TL_12_3;
wire wire_in_cluster_sb_TL_12_4;
wire wire_in_cluster_sb_TL_12_5;
wire wire_in_cluster_sb_TL_12_6;
wire wire_in_cluster_sb_TL_12_7;
wire wire_in_cluster_sb_TL_12_8;
wire wire_in_cluster_sb_TL_12_9;
wire wire_in_cluster_sb_TL_13_0;
wire wire_in_cluster_sb_TL_13_1;
wire wire_in_cluster_sb_TL_13_10;
wire wire_in_cluster_sb_TL_13_11;
wire wire_in_cluster_sb_TL_13_12;
wire wire_in_cluster_sb_TL_13_13;
wire wire_in_cluster_sb_TL_13_14;
wire wire_in_cluster_sb_TL_13_15;
wire wire_in_cluster_sb_TL_13_2;
wire wire_in_cluster_sb_TL_13_3;
wire wire_in_cluster_sb_TL_13_4;
wire wire_in_cluster_sb_TL_13_5;
wire wire_in_cluster_sb_TL_13_6;
wire wire_in_cluster_sb_TL_13_7;
wire wire_in_cluster_sb_TL_13_8;
wire wire_in_cluster_sb_TL_13_9;
wire wire_in_cluster_sb_TL_14_0;
wire wire_in_cluster_sb_TL_14_1;
wire wire_in_cluster_sb_TL_14_10;
wire wire_in_cluster_sb_TL_14_11;
wire wire_in_cluster_sb_TL_14_12;
wire wire_in_cluster_sb_TL_14_13;
wire wire_in_cluster_sb_TL_14_14;
wire wire_in_cluster_sb_TL_14_15;
wire wire_in_cluster_sb_TL_14_2;
wire wire_in_cluster_sb_TL_14_3;
wire wire_in_cluster_sb_TL_14_4;
wire wire_in_cluster_sb_TL_14_5;
wire wire_in_cluster_sb_TL_14_6;
wire wire_in_cluster_sb_TL_14_7;
wire wire_in_cluster_sb_TL_14_8;
wire wire_in_cluster_sb_TL_14_9;
wire wire_in_cluster_sb_TL_15_0;
wire wire_in_cluster_sb_TL_15_1;
wire wire_in_cluster_sb_TL_15_10;
wire wire_in_cluster_sb_TL_15_11;
wire wire_in_cluster_sb_TL_15_12;
wire wire_in_cluster_sb_TL_15_13;
wire wire_in_cluster_sb_TL_15_14;
wire wire_in_cluster_sb_TL_15_15;
wire wire_in_cluster_sb_TL_15_2;
wire wire_in_cluster_sb_TL_15_3;
wire wire_in_cluster_sb_TL_15_4;
wire wire_in_cluster_sb_TL_15_5;
wire wire_in_cluster_sb_TL_15_6;
wire wire_in_cluster_sb_TL_15_7;
wire wire_in_cluster_sb_TL_15_8;
wire wire_in_cluster_sb_TL_15_9;
wire wire_in_cluster_sb_TL_1_0;
wire wire_in_cluster_sb_TL_1_1;
wire wire_in_cluster_sb_TL_1_10;
wire wire_in_cluster_sb_TL_1_11;
wire wire_in_cluster_sb_TL_1_12;
wire wire_in_cluster_sb_TL_1_13;
wire wire_in_cluster_sb_TL_1_14;
wire wire_in_cluster_sb_TL_1_15;
wire wire_in_cluster_sb_TL_1_2;
wire wire_in_cluster_sb_TL_1_3;
wire wire_in_cluster_sb_TL_1_4;
wire wire_in_cluster_sb_TL_1_5;
wire wire_in_cluster_sb_TL_1_6;
wire wire_in_cluster_sb_TL_1_7;
wire wire_in_cluster_sb_TL_1_8;
wire wire_in_cluster_sb_TL_1_9;
wire wire_in_cluster_sb_TL_2_0;
wire wire_in_cluster_sb_TL_2_1;
wire wire_in_cluster_sb_TL_2_10;
wire wire_in_cluster_sb_TL_2_11;
wire wire_in_cluster_sb_TL_2_12;
wire wire_in_cluster_sb_TL_2_13;
wire wire_in_cluster_sb_TL_2_14;
wire wire_in_cluster_sb_TL_2_15;
wire wire_in_cluster_sb_TL_2_2;
wire wire_in_cluster_sb_TL_2_3;
wire wire_in_cluster_sb_TL_2_4;
wire wire_in_cluster_sb_TL_2_5;
wire wire_in_cluster_sb_TL_2_6;
wire wire_in_cluster_sb_TL_2_7;
wire wire_in_cluster_sb_TL_2_8;
wire wire_in_cluster_sb_TL_2_9;
wire wire_in_cluster_sb_TL_3_0;
wire wire_in_cluster_sb_TL_3_1;
wire wire_in_cluster_sb_TL_3_10;
wire wire_in_cluster_sb_TL_3_11;
wire wire_in_cluster_sb_TL_3_12;
wire wire_in_cluster_sb_TL_3_13;
wire wire_in_cluster_sb_TL_3_14;
wire wire_in_cluster_sb_TL_3_15;
wire wire_in_cluster_sb_TL_3_2;
wire wire_in_cluster_sb_TL_3_3;
wire wire_in_cluster_sb_TL_3_4;
wire wire_in_cluster_sb_TL_3_5;
wire wire_in_cluster_sb_TL_3_6;
wire wire_in_cluster_sb_TL_3_7;
wire wire_in_cluster_sb_TL_3_8;
wire wire_in_cluster_sb_TL_3_9;
wire wire_in_cluster_sb_TL_4_0;
wire wire_in_cluster_sb_TL_4_1;
wire wire_in_cluster_sb_TL_4_10;
wire wire_in_cluster_sb_TL_4_11;
wire wire_in_cluster_sb_TL_4_12;
wire wire_in_cluster_sb_TL_4_13;
wire wire_in_cluster_sb_TL_4_14;
wire wire_in_cluster_sb_TL_4_15;
wire wire_in_cluster_sb_TL_4_2;
wire wire_in_cluster_sb_TL_4_3;
wire wire_in_cluster_sb_TL_4_4;
wire wire_in_cluster_sb_TL_4_5;
wire wire_in_cluster_sb_TL_4_6;
wire wire_in_cluster_sb_TL_4_7;
wire wire_in_cluster_sb_TL_4_8;
wire wire_in_cluster_sb_TL_4_9;
wire wire_in_cluster_sb_TL_5_0;
wire wire_in_cluster_sb_TL_5_1;
wire wire_in_cluster_sb_TL_5_10;
wire wire_in_cluster_sb_TL_5_11;
wire wire_in_cluster_sb_TL_5_12;
wire wire_in_cluster_sb_TL_5_13;
wire wire_in_cluster_sb_TL_5_14;
wire wire_in_cluster_sb_TL_5_15;
wire wire_in_cluster_sb_TL_5_2;
wire wire_in_cluster_sb_TL_5_3;
wire wire_in_cluster_sb_TL_5_4;
wire wire_in_cluster_sb_TL_5_5;
wire wire_in_cluster_sb_TL_5_6;
wire wire_in_cluster_sb_TL_5_7;
wire wire_in_cluster_sb_TL_5_8;
wire wire_in_cluster_sb_TL_5_9;
wire wire_in_cluster_sb_TL_6_0;
wire wire_in_cluster_sb_TL_6_1;
wire wire_in_cluster_sb_TL_6_10;
wire wire_in_cluster_sb_TL_6_11;
wire wire_in_cluster_sb_TL_6_12;
wire wire_in_cluster_sb_TL_6_13;
wire wire_in_cluster_sb_TL_6_14;
wire wire_in_cluster_sb_TL_6_15;
wire wire_in_cluster_sb_TL_6_2;
wire wire_in_cluster_sb_TL_6_3;
wire wire_in_cluster_sb_TL_6_4;
wire wire_in_cluster_sb_TL_6_5;
wire wire_in_cluster_sb_TL_6_6;
wire wire_in_cluster_sb_TL_6_7;
wire wire_in_cluster_sb_TL_6_8;
wire wire_in_cluster_sb_TL_6_9;
wire wire_in_cluster_sb_TL_7_0;
wire wire_in_cluster_sb_TL_7_1;
wire wire_in_cluster_sb_TL_7_10;
wire wire_in_cluster_sb_TL_7_11;
wire wire_in_cluster_sb_TL_7_12;
wire wire_in_cluster_sb_TL_7_13;
wire wire_in_cluster_sb_TL_7_14;
wire wire_in_cluster_sb_TL_7_15;
wire wire_in_cluster_sb_TL_7_2;
wire wire_in_cluster_sb_TL_7_3;
wire wire_in_cluster_sb_TL_7_4;
wire wire_in_cluster_sb_TL_7_5;
wire wire_in_cluster_sb_TL_7_6;
wire wire_in_cluster_sb_TL_7_7;
wire wire_in_cluster_sb_TL_7_8;
wire wire_in_cluster_sb_TL_7_9;
wire wire_in_cluster_sb_TL_8_0;
wire wire_in_cluster_sb_TL_8_1;
wire wire_in_cluster_sb_TL_8_10;
wire wire_in_cluster_sb_TL_8_11;
wire wire_in_cluster_sb_TL_8_12;
wire wire_in_cluster_sb_TL_8_13;
wire wire_in_cluster_sb_TL_8_14;
wire wire_in_cluster_sb_TL_8_15;
wire wire_in_cluster_sb_TL_8_2;
wire wire_in_cluster_sb_TL_8_3;
wire wire_in_cluster_sb_TL_8_4;
wire wire_in_cluster_sb_TL_8_5;
wire wire_in_cluster_sb_TL_8_6;
wire wire_in_cluster_sb_TL_8_7;
wire wire_in_cluster_sb_TL_8_8;
wire wire_in_cluster_sb_TL_8_9;
wire wire_in_cluster_sb_TL_9_0;
wire wire_in_cluster_sb_TL_9_1;
wire wire_in_cluster_sb_TL_9_10;
wire wire_in_cluster_sb_TL_9_11;
wire wire_in_cluster_sb_TL_9_12;
wire wire_in_cluster_sb_TL_9_13;
wire wire_in_cluster_sb_TL_9_14;
wire wire_in_cluster_sb_TL_9_15;
wire wire_in_cluster_sb_TL_9_2;
wire wire_in_cluster_sb_TL_9_3;
wire wire_in_cluster_sb_TL_9_4;
wire wire_in_cluster_sb_TL_9_5;
wire wire_in_cluster_sb_TL_9_6;
wire wire_in_cluster_sb_TL_9_7;
wire wire_in_cluster_sb_TL_9_8;
wire wire_in_cluster_sb_TL_9_9;
wire wire_out_cluster_sb_BL_0_0;
wire wire_out_cluster_sb_BL_0_1;
wire wire_out_cluster_sb_BL_0_10;
wire wire_out_cluster_sb_BL_0_11;
wire wire_out_cluster_sb_BL_0_12;
wire wire_out_cluster_sb_BL_0_13;
wire wire_out_cluster_sb_BL_0_14;
wire wire_out_cluster_sb_BL_0_15;
wire wire_out_cluster_sb_BL_0_2;
wire wire_out_cluster_sb_BL_0_3;
wire wire_out_cluster_sb_BL_0_4;
wire wire_out_cluster_sb_BL_0_5;
wire wire_out_cluster_sb_BL_0_6;
wire wire_out_cluster_sb_BL_0_7;
wire wire_out_cluster_sb_BL_0_8;
wire wire_out_cluster_sb_BL_0_9;
wire wire_out_cluster_sb_BL_1_0;
wire wire_out_cluster_sb_BL_1_1;
wire wire_out_cluster_sb_BL_1_10;
wire wire_out_cluster_sb_BL_1_11;
wire wire_out_cluster_sb_BL_1_12;
wire wire_out_cluster_sb_BL_1_13;
wire wire_out_cluster_sb_BL_1_14;
wire wire_out_cluster_sb_BL_1_15;
wire wire_out_cluster_sb_BL_1_2;
wire wire_out_cluster_sb_BL_1_3;
wire wire_out_cluster_sb_BL_1_4;
wire wire_out_cluster_sb_BL_1_5;
wire wire_out_cluster_sb_BL_1_6;
wire wire_out_cluster_sb_BL_1_7;
wire wire_out_cluster_sb_BL_1_8;
wire wire_out_cluster_sb_BL_1_9;
wire wire_out_cluster_sb_BL_2_0;
wire wire_out_cluster_sb_BL_2_1;
wire wire_out_cluster_sb_BL_2_10;
wire wire_out_cluster_sb_BL_2_11;
wire wire_out_cluster_sb_BL_2_12;
wire wire_out_cluster_sb_BL_2_13;
wire wire_out_cluster_sb_BL_2_14;
wire wire_out_cluster_sb_BL_2_15;
wire wire_out_cluster_sb_BL_2_2;
wire wire_out_cluster_sb_BL_2_3;
wire wire_out_cluster_sb_BL_2_4;
wire wire_out_cluster_sb_BL_2_5;
wire wire_out_cluster_sb_BL_2_6;
wire wire_out_cluster_sb_BL_2_7;
wire wire_out_cluster_sb_BL_2_8;
wire wire_out_cluster_sb_BL_2_9;
wire wire_out_cluster_sb_BL_3_0;
wire wire_out_cluster_sb_BL_3_1;
wire wire_out_cluster_sb_BL_3_10;
wire wire_out_cluster_sb_BL_3_11;
wire wire_out_cluster_sb_BL_3_12;
wire wire_out_cluster_sb_BL_3_13;
wire wire_out_cluster_sb_BL_3_14;
wire wire_out_cluster_sb_BL_3_15;
wire wire_out_cluster_sb_BL_3_2;
wire wire_out_cluster_sb_BL_3_3;
wire wire_out_cluster_sb_BL_3_4;
wire wire_out_cluster_sb_BL_3_5;
wire wire_out_cluster_sb_BL_3_6;
wire wire_out_cluster_sb_BL_3_7;
wire wire_out_cluster_sb_BL_3_8;
wire wire_out_cluster_sb_BL_3_9;
wire wire_out_cluster_sb_BR_0_0;
wire wire_out_cluster_sb_BR_0_1;
wire wire_out_cluster_sb_BR_0_10;
wire wire_out_cluster_sb_BR_0_11;
wire wire_out_cluster_sb_BR_0_12;
wire wire_out_cluster_sb_BR_0_13;
wire wire_out_cluster_sb_BR_0_14;
wire wire_out_cluster_sb_BR_0_15;
wire wire_out_cluster_sb_BR_0_2;
wire wire_out_cluster_sb_BR_0_3;
wire wire_out_cluster_sb_BR_0_4;
wire wire_out_cluster_sb_BR_0_5;
wire wire_out_cluster_sb_BR_0_6;
wire wire_out_cluster_sb_BR_0_7;
wire wire_out_cluster_sb_BR_0_8;
wire wire_out_cluster_sb_BR_0_9;
wire wire_out_cluster_sb_BR_1_0;
wire wire_out_cluster_sb_BR_1_1;
wire wire_out_cluster_sb_BR_1_10;
wire wire_out_cluster_sb_BR_1_11;
wire wire_out_cluster_sb_BR_1_12;
wire wire_out_cluster_sb_BR_1_13;
wire wire_out_cluster_sb_BR_1_14;
wire wire_out_cluster_sb_BR_1_15;
wire wire_out_cluster_sb_BR_1_2;
wire wire_out_cluster_sb_BR_1_3;
wire wire_out_cluster_sb_BR_1_4;
wire wire_out_cluster_sb_BR_1_5;
wire wire_out_cluster_sb_BR_1_6;
wire wire_out_cluster_sb_BR_1_7;
wire wire_out_cluster_sb_BR_1_8;
wire wire_out_cluster_sb_BR_1_9;
wire wire_out_cluster_sb_BR_2_0;
wire wire_out_cluster_sb_BR_2_1;
wire wire_out_cluster_sb_BR_2_10;
wire wire_out_cluster_sb_BR_2_11;
wire wire_out_cluster_sb_BR_2_12;
wire wire_out_cluster_sb_BR_2_13;
wire wire_out_cluster_sb_BR_2_14;
wire wire_out_cluster_sb_BR_2_15;
wire wire_out_cluster_sb_BR_2_2;
wire wire_out_cluster_sb_BR_2_3;
wire wire_out_cluster_sb_BR_2_4;
wire wire_out_cluster_sb_BR_2_5;
wire wire_out_cluster_sb_BR_2_6;
wire wire_out_cluster_sb_BR_2_7;
wire wire_out_cluster_sb_BR_2_8;
wire wire_out_cluster_sb_BR_2_9;
wire wire_out_cluster_sb_BR_3_0;
wire wire_out_cluster_sb_BR_3_1;
wire wire_out_cluster_sb_BR_3_10;
wire wire_out_cluster_sb_BR_3_11;
wire wire_out_cluster_sb_BR_3_12;
wire wire_out_cluster_sb_BR_3_13;
wire wire_out_cluster_sb_BR_3_14;
wire wire_out_cluster_sb_BR_3_15;
wire wire_out_cluster_sb_BR_3_2;
wire wire_out_cluster_sb_BR_3_3;
wire wire_out_cluster_sb_BR_3_4;
wire wire_out_cluster_sb_BR_3_5;
wire wire_out_cluster_sb_BR_3_6;
wire wire_out_cluster_sb_BR_3_7;
wire wire_out_cluster_sb_BR_3_8;
wire wire_out_cluster_sb_BR_3_9;
wire wire_out_cluster_sb_TL_0_0;
wire wire_out_cluster_sb_TL_0_1;
wire wire_out_cluster_sb_TL_0_10;
wire wire_out_cluster_sb_TL_0_11;
wire wire_out_cluster_sb_TL_0_12;
wire wire_out_cluster_sb_TL_0_13;
wire wire_out_cluster_sb_TL_0_14;
wire wire_out_cluster_sb_TL_0_15;
wire wire_out_cluster_sb_TL_0_2;
wire wire_out_cluster_sb_TL_0_3;
wire wire_out_cluster_sb_TL_0_4;
wire wire_out_cluster_sb_TL_0_5;
wire wire_out_cluster_sb_TL_0_6;
wire wire_out_cluster_sb_TL_0_7;
wire wire_out_cluster_sb_TL_0_8;
wire wire_out_cluster_sb_TL_0_9;
wire wire_out_cluster_sb_TL_1_0;
wire wire_out_cluster_sb_TL_1_1;
wire wire_out_cluster_sb_TL_1_10;
wire wire_out_cluster_sb_TL_1_11;
wire wire_out_cluster_sb_TL_1_12;
wire wire_out_cluster_sb_TL_1_13;
wire wire_out_cluster_sb_TL_1_14;
wire wire_out_cluster_sb_TL_1_15;
wire wire_out_cluster_sb_TL_1_2;
wire wire_out_cluster_sb_TL_1_3;
wire wire_out_cluster_sb_TL_1_4;
wire wire_out_cluster_sb_TL_1_5;
wire wire_out_cluster_sb_TL_1_6;
wire wire_out_cluster_sb_TL_1_7;
wire wire_out_cluster_sb_TL_1_8;
wire wire_out_cluster_sb_TL_1_9;
wire wire_out_cluster_sb_TL_2_0;
wire wire_out_cluster_sb_TL_2_1;
wire wire_out_cluster_sb_TL_2_10;
wire wire_out_cluster_sb_TL_2_11;
wire wire_out_cluster_sb_TL_2_12;
wire wire_out_cluster_sb_TL_2_13;
wire wire_out_cluster_sb_TL_2_14;
wire wire_out_cluster_sb_TL_2_15;
wire wire_out_cluster_sb_TL_2_2;
wire wire_out_cluster_sb_TL_2_3;
wire wire_out_cluster_sb_TL_2_4;
wire wire_out_cluster_sb_TL_2_5;
wire wire_out_cluster_sb_TL_2_6;
wire wire_out_cluster_sb_TL_2_7;
wire wire_out_cluster_sb_TL_2_8;
wire wire_out_cluster_sb_TL_2_9;
wire wire_out_cluster_sb_TL_3_0;
wire wire_out_cluster_sb_TL_3_1;
wire wire_out_cluster_sb_TL_3_10;
wire wire_out_cluster_sb_TL_3_11;
wire wire_out_cluster_sb_TL_3_12;
wire wire_out_cluster_sb_TL_3_13;
wire wire_out_cluster_sb_TL_3_14;
wire wire_out_cluster_sb_TL_3_15;
wire wire_out_cluster_sb_TL_3_2;
wire wire_out_cluster_sb_TL_3_3;
wire wire_out_cluster_sb_TL_3_4;
wire wire_out_cluster_sb_TL_3_5;
wire wire_out_cluster_sb_TL_3_6;
wire wire_out_cluster_sb_TL_3_7;
wire wire_out_cluster_sb_TL_3_8;
wire wire_out_cluster_sb_TL_3_9;
wire wire_sb_bottom_input_0_0;
wire wire_sb_bottom_input_0_1;
wire wire_sb_bottom_input_0_10;
wire wire_sb_bottom_input_0_11;
wire wire_sb_bottom_input_0_12;
wire wire_sb_bottom_input_0_13;
wire wire_sb_bottom_input_0_14;
wire wire_sb_bottom_input_0_15;
wire wire_sb_bottom_input_0_16;
wire wire_sb_bottom_input_0_17;
wire wire_sb_bottom_input_0_18;
wire wire_sb_bottom_input_0_19;
wire wire_sb_bottom_input_0_2;
wire wire_sb_bottom_input_0_3;
wire wire_sb_bottom_input_0_4;
wire wire_sb_bottom_input_0_5;
wire wire_sb_bottom_input_0_6;
wire wire_sb_bottom_input_0_7;
wire wire_sb_bottom_input_0_8;
wire wire_sb_bottom_input_0_9;
wire wire_sb_bottom_input_10_0;
wire wire_sb_bottom_input_10_1;
wire wire_sb_bottom_input_10_10;
wire wire_sb_bottom_input_10_11;
wire wire_sb_bottom_input_10_12;
wire wire_sb_bottom_input_10_13;
wire wire_sb_bottom_input_10_14;
wire wire_sb_bottom_input_10_15;
wire wire_sb_bottom_input_10_16;
wire wire_sb_bottom_input_10_17;
wire wire_sb_bottom_input_10_18;
wire wire_sb_bottom_input_10_19;
wire wire_sb_bottom_input_10_2;
wire wire_sb_bottom_input_10_3;
wire wire_sb_bottom_input_10_4;
wire wire_sb_bottom_input_10_5;
wire wire_sb_bottom_input_10_6;
wire wire_sb_bottom_input_10_7;
wire wire_sb_bottom_input_10_8;
wire wire_sb_bottom_input_10_9;
wire wire_sb_bottom_input_11_0;
wire wire_sb_bottom_input_11_1;
wire wire_sb_bottom_input_11_10;
wire wire_sb_bottom_input_11_11;
wire wire_sb_bottom_input_11_12;
wire wire_sb_bottom_input_11_13;
wire wire_sb_bottom_input_11_14;
wire wire_sb_bottom_input_11_15;
wire wire_sb_bottom_input_11_16;
wire wire_sb_bottom_input_11_17;
wire wire_sb_bottom_input_11_18;
wire wire_sb_bottom_input_11_19;
wire wire_sb_bottom_input_11_2;
wire wire_sb_bottom_input_11_3;
wire wire_sb_bottom_input_11_4;
wire wire_sb_bottom_input_11_5;
wire wire_sb_bottom_input_11_6;
wire wire_sb_bottom_input_11_7;
wire wire_sb_bottom_input_11_8;
wire wire_sb_bottom_input_11_9;
wire wire_sb_bottom_input_1_0;
wire wire_sb_bottom_input_1_1;
wire wire_sb_bottom_input_1_10;
wire wire_sb_bottom_input_1_11;
wire wire_sb_bottom_input_1_12;
wire wire_sb_bottom_input_1_13;
wire wire_sb_bottom_input_1_14;
wire wire_sb_bottom_input_1_15;
wire wire_sb_bottom_input_1_16;
wire wire_sb_bottom_input_1_17;
wire wire_sb_bottom_input_1_18;
wire wire_sb_bottom_input_1_19;
wire wire_sb_bottom_input_1_2;
wire wire_sb_bottom_input_1_3;
wire wire_sb_bottom_input_1_4;
wire wire_sb_bottom_input_1_5;
wire wire_sb_bottom_input_1_6;
wire wire_sb_bottom_input_1_7;
wire wire_sb_bottom_input_1_8;
wire wire_sb_bottom_input_1_9;
wire wire_sb_bottom_input_2_0;
wire wire_sb_bottom_input_2_1;
wire wire_sb_bottom_input_2_10;
wire wire_sb_bottom_input_2_11;
wire wire_sb_bottom_input_2_12;
wire wire_sb_bottom_input_2_13;
wire wire_sb_bottom_input_2_14;
wire wire_sb_bottom_input_2_15;
wire wire_sb_bottom_input_2_16;
wire wire_sb_bottom_input_2_17;
wire wire_sb_bottom_input_2_18;
wire wire_sb_bottom_input_2_19;
wire wire_sb_bottom_input_2_2;
wire wire_sb_bottom_input_2_3;
wire wire_sb_bottom_input_2_4;
wire wire_sb_bottom_input_2_5;
wire wire_sb_bottom_input_2_6;
wire wire_sb_bottom_input_2_7;
wire wire_sb_bottom_input_2_8;
wire wire_sb_bottom_input_2_9;
wire wire_sb_bottom_input_3_0;
wire wire_sb_bottom_input_3_1;
wire wire_sb_bottom_input_3_10;
wire wire_sb_bottom_input_3_11;
wire wire_sb_bottom_input_3_12;
wire wire_sb_bottom_input_3_13;
wire wire_sb_bottom_input_3_14;
wire wire_sb_bottom_input_3_15;
wire wire_sb_bottom_input_3_16;
wire wire_sb_bottom_input_3_17;
wire wire_sb_bottom_input_3_18;
wire wire_sb_bottom_input_3_19;
wire wire_sb_bottom_input_3_2;
wire wire_sb_bottom_input_3_3;
wire wire_sb_bottom_input_3_4;
wire wire_sb_bottom_input_3_5;
wire wire_sb_bottom_input_3_6;
wire wire_sb_bottom_input_3_7;
wire wire_sb_bottom_input_3_8;
wire wire_sb_bottom_input_3_9;
wire wire_sb_bottom_input_4_0;
wire wire_sb_bottom_input_4_1;
wire wire_sb_bottom_input_4_10;
wire wire_sb_bottom_input_4_11;
wire wire_sb_bottom_input_4_12;
wire wire_sb_bottom_input_4_13;
wire wire_sb_bottom_input_4_14;
wire wire_sb_bottom_input_4_15;
wire wire_sb_bottom_input_4_16;
wire wire_sb_bottom_input_4_17;
wire wire_sb_bottom_input_4_18;
wire wire_sb_bottom_input_4_19;
wire wire_sb_bottom_input_4_2;
wire wire_sb_bottom_input_4_3;
wire wire_sb_bottom_input_4_4;
wire wire_sb_bottom_input_4_5;
wire wire_sb_bottom_input_4_6;
wire wire_sb_bottom_input_4_7;
wire wire_sb_bottom_input_4_8;
wire wire_sb_bottom_input_4_9;
wire wire_sb_bottom_input_5_0;
wire wire_sb_bottom_input_5_1;
wire wire_sb_bottom_input_5_10;
wire wire_sb_bottom_input_5_11;
wire wire_sb_bottom_input_5_12;
wire wire_sb_bottom_input_5_13;
wire wire_sb_bottom_input_5_14;
wire wire_sb_bottom_input_5_15;
wire wire_sb_bottom_input_5_16;
wire wire_sb_bottom_input_5_17;
wire wire_sb_bottom_input_5_18;
wire wire_sb_bottom_input_5_19;
wire wire_sb_bottom_input_5_2;
wire wire_sb_bottom_input_5_3;
wire wire_sb_bottom_input_5_4;
wire wire_sb_bottom_input_5_5;
wire wire_sb_bottom_input_5_6;
wire wire_sb_bottom_input_5_7;
wire wire_sb_bottom_input_5_8;
wire wire_sb_bottom_input_5_9;
wire wire_sb_bottom_input_6_0;
wire wire_sb_bottom_input_6_1;
wire wire_sb_bottom_input_6_10;
wire wire_sb_bottom_input_6_11;
wire wire_sb_bottom_input_6_12;
wire wire_sb_bottom_input_6_13;
wire wire_sb_bottom_input_6_14;
wire wire_sb_bottom_input_6_15;
wire wire_sb_bottom_input_6_16;
wire wire_sb_bottom_input_6_17;
wire wire_sb_bottom_input_6_18;
wire wire_sb_bottom_input_6_19;
wire wire_sb_bottom_input_6_2;
wire wire_sb_bottom_input_6_3;
wire wire_sb_bottom_input_6_4;
wire wire_sb_bottom_input_6_5;
wire wire_sb_bottom_input_6_6;
wire wire_sb_bottom_input_6_7;
wire wire_sb_bottom_input_6_8;
wire wire_sb_bottom_input_6_9;
wire wire_sb_bottom_input_7_0;
wire wire_sb_bottom_input_7_1;
wire wire_sb_bottom_input_7_10;
wire wire_sb_bottom_input_7_11;
wire wire_sb_bottom_input_7_12;
wire wire_sb_bottom_input_7_13;
wire wire_sb_bottom_input_7_14;
wire wire_sb_bottom_input_7_15;
wire wire_sb_bottom_input_7_16;
wire wire_sb_bottom_input_7_17;
wire wire_sb_bottom_input_7_18;
wire wire_sb_bottom_input_7_19;
wire wire_sb_bottom_input_7_2;
wire wire_sb_bottom_input_7_3;
wire wire_sb_bottom_input_7_4;
wire wire_sb_bottom_input_7_5;
wire wire_sb_bottom_input_7_6;
wire wire_sb_bottom_input_7_7;
wire wire_sb_bottom_input_7_8;
wire wire_sb_bottom_input_7_9;
wire wire_sb_bottom_input_8_0;
wire wire_sb_bottom_input_8_1;
wire wire_sb_bottom_input_8_10;
wire wire_sb_bottom_input_8_11;
wire wire_sb_bottom_input_8_12;
wire wire_sb_bottom_input_8_13;
wire wire_sb_bottom_input_8_14;
wire wire_sb_bottom_input_8_15;
wire wire_sb_bottom_input_8_16;
wire wire_sb_bottom_input_8_17;
wire wire_sb_bottom_input_8_18;
wire wire_sb_bottom_input_8_19;
wire wire_sb_bottom_input_8_2;
wire wire_sb_bottom_input_8_3;
wire wire_sb_bottom_input_8_4;
wire wire_sb_bottom_input_8_5;
wire wire_sb_bottom_input_8_6;
wire wire_sb_bottom_input_8_7;
wire wire_sb_bottom_input_8_8;
wire wire_sb_bottom_input_8_9;
wire wire_sb_bottom_input_9_0;
wire wire_sb_bottom_input_9_1;
wire wire_sb_bottom_input_9_10;
wire wire_sb_bottom_input_9_11;
wire wire_sb_bottom_input_9_12;
wire wire_sb_bottom_input_9_13;
wire wire_sb_bottom_input_9_14;
wire wire_sb_bottom_input_9_15;
wire wire_sb_bottom_input_9_16;
wire wire_sb_bottom_input_9_17;
wire wire_sb_bottom_input_9_18;
wire wire_sb_bottom_input_9_19;
wire wire_sb_bottom_input_9_2;
wire wire_sb_bottom_input_9_3;
wire wire_sb_bottom_input_9_4;
wire wire_sb_bottom_input_9_5;
wire wire_sb_bottom_input_9_6;
wire wire_sb_bottom_input_9_7;
wire wire_sb_bottom_input_9_8;
wire wire_sb_bottom_input_9_9;
wire wire_sb_bottom_output_0_0;
wire wire_sb_bottom_output_0_1;
wire wire_sb_bottom_output_0_10;
wire wire_sb_bottom_output_0_11;
wire wire_sb_bottom_output_0_12;
wire wire_sb_bottom_output_0_13;
wire wire_sb_bottom_output_0_14;
wire wire_sb_bottom_output_0_15;
wire wire_sb_bottom_output_0_16;
wire wire_sb_bottom_output_0_17;
wire wire_sb_bottom_output_0_18;
wire wire_sb_bottom_output_0_19;
wire wire_sb_bottom_output_0_2;
wire wire_sb_bottom_output_0_3;
wire wire_sb_bottom_output_0_4;
wire wire_sb_bottom_output_0_5;
wire wire_sb_bottom_output_0_6;
wire wire_sb_bottom_output_0_7;
wire wire_sb_bottom_output_0_8;
wire wire_sb_bottom_output_0_9;
wire wire_sb_bottom_output_10_0;
wire wire_sb_bottom_output_10_1;
wire wire_sb_bottom_output_10_10;
wire wire_sb_bottom_output_10_11;
wire wire_sb_bottom_output_10_12;
wire wire_sb_bottom_output_10_13;
wire wire_sb_bottom_output_10_14;
wire wire_sb_bottom_output_10_15;
wire wire_sb_bottom_output_10_16;
wire wire_sb_bottom_output_10_17;
wire wire_sb_bottom_output_10_18;
wire wire_sb_bottom_output_10_19;
wire wire_sb_bottom_output_10_2;
wire wire_sb_bottom_output_10_3;
wire wire_sb_bottom_output_10_4;
wire wire_sb_bottom_output_10_5;
wire wire_sb_bottom_output_10_6;
wire wire_sb_bottom_output_10_7;
wire wire_sb_bottom_output_10_8;
wire wire_sb_bottom_output_10_9;
wire wire_sb_bottom_output_11_0;
wire wire_sb_bottom_output_11_1;
wire wire_sb_bottom_output_11_10;
wire wire_sb_bottom_output_11_11;
wire wire_sb_bottom_output_11_12;
wire wire_sb_bottom_output_11_13;
wire wire_sb_bottom_output_11_14;
wire wire_sb_bottom_output_11_15;
wire wire_sb_bottom_output_11_16;
wire wire_sb_bottom_output_11_17;
wire wire_sb_bottom_output_11_18;
wire wire_sb_bottom_output_11_19;
wire wire_sb_bottom_output_11_2;
wire wire_sb_bottom_output_11_3;
wire wire_sb_bottom_output_11_4;
wire wire_sb_bottom_output_11_5;
wire wire_sb_bottom_output_11_6;
wire wire_sb_bottom_output_11_7;
wire wire_sb_bottom_output_11_8;
wire wire_sb_bottom_output_11_9;
wire wire_sb_bottom_output_1_0;
wire wire_sb_bottom_output_1_1;
wire wire_sb_bottom_output_1_10;
wire wire_sb_bottom_output_1_11;
wire wire_sb_bottom_output_1_12;
wire wire_sb_bottom_output_1_13;
wire wire_sb_bottom_output_1_14;
wire wire_sb_bottom_output_1_15;
wire wire_sb_bottom_output_1_16;
wire wire_sb_bottom_output_1_17;
wire wire_sb_bottom_output_1_18;
wire wire_sb_bottom_output_1_19;
wire wire_sb_bottom_output_1_2;
wire wire_sb_bottom_output_1_3;
wire wire_sb_bottom_output_1_4;
wire wire_sb_bottom_output_1_5;
wire wire_sb_bottom_output_1_6;
wire wire_sb_bottom_output_1_7;
wire wire_sb_bottom_output_1_8;
wire wire_sb_bottom_output_1_9;
wire wire_sb_bottom_output_2_0;
wire wire_sb_bottom_output_2_1;
wire wire_sb_bottom_output_2_10;
wire wire_sb_bottom_output_2_11;
wire wire_sb_bottom_output_2_12;
wire wire_sb_bottom_output_2_13;
wire wire_sb_bottom_output_2_14;
wire wire_sb_bottom_output_2_15;
wire wire_sb_bottom_output_2_16;
wire wire_sb_bottom_output_2_17;
wire wire_sb_bottom_output_2_18;
wire wire_sb_bottom_output_2_19;
wire wire_sb_bottom_output_2_2;
wire wire_sb_bottom_output_2_3;
wire wire_sb_bottom_output_2_4;
wire wire_sb_bottom_output_2_5;
wire wire_sb_bottom_output_2_6;
wire wire_sb_bottom_output_2_7;
wire wire_sb_bottom_output_2_8;
wire wire_sb_bottom_output_2_9;
wire wire_sb_bottom_output_3_0;
wire wire_sb_bottom_output_3_1;
wire wire_sb_bottom_output_3_10;
wire wire_sb_bottom_output_3_11;
wire wire_sb_bottom_output_3_12;
wire wire_sb_bottom_output_3_13;
wire wire_sb_bottom_output_3_14;
wire wire_sb_bottom_output_3_15;
wire wire_sb_bottom_output_3_16;
wire wire_sb_bottom_output_3_17;
wire wire_sb_bottom_output_3_18;
wire wire_sb_bottom_output_3_19;
wire wire_sb_bottom_output_3_2;
wire wire_sb_bottom_output_3_3;
wire wire_sb_bottom_output_3_4;
wire wire_sb_bottom_output_3_5;
wire wire_sb_bottom_output_3_6;
wire wire_sb_bottom_output_3_7;
wire wire_sb_bottom_output_3_8;
wire wire_sb_bottom_output_3_9;
wire wire_sb_bottom_output_4_0;
wire wire_sb_bottom_output_4_1;
wire wire_sb_bottom_output_4_10;
wire wire_sb_bottom_output_4_11;
wire wire_sb_bottom_output_4_12;
wire wire_sb_bottom_output_4_13;
wire wire_sb_bottom_output_4_14;
wire wire_sb_bottom_output_4_15;
wire wire_sb_bottom_output_4_16;
wire wire_sb_bottom_output_4_17;
wire wire_sb_bottom_output_4_18;
wire wire_sb_bottom_output_4_19;
wire wire_sb_bottom_output_4_2;
wire wire_sb_bottom_output_4_3;
wire wire_sb_bottom_output_4_4;
wire wire_sb_bottom_output_4_5;
wire wire_sb_bottom_output_4_6;
wire wire_sb_bottom_output_4_7;
wire wire_sb_bottom_output_4_8;
wire wire_sb_bottom_output_4_9;
wire wire_sb_bottom_output_5_0;
wire wire_sb_bottom_output_5_1;
wire wire_sb_bottom_output_5_10;
wire wire_sb_bottom_output_5_11;
wire wire_sb_bottom_output_5_12;
wire wire_sb_bottom_output_5_13;
wire wire_sb_bottom_output_5_14;
wire wire_sb_bottom_output_5_15;
wire wire_sb_bottom_output_5_16;
wire wire_sb_bottom_output_5_17;
wire wire_sb_bottom_output_5_18;
wire wire_sb_bottom_output_5_19;
wire wire_sb_bottom_output_5_2;
wire wire_sb_bottom_output_5_3;
wire wire_sb_bottom_output_5_4;
wire wire_sb_bottom_output_5_5;
wire wire_sb_bottom_output_5_6;
wire wire_sb_bottom_output_5_7;
wire wire_sb_bottom_output_5_8;
wire wire_sb_bottom_output_5_9;
wire wire_sb_bottom_output_6_0;
wire wire_sb_bottom_output_6_1;
wire wire_sb_bottom_output_6_10;
wire wire_sb_bottom_output_6_11;
wire wire_sb_bottom_output_6_12;
wire wire_sb_bottom_output_6_13;
wire wire_sb_bottom_output_6_14;
wire wire_sb_bottom_output_6_15;
wire wire_sb_bottom_output_6_16;
wire wire_sb_bottom_output_6_17;
wire wire_sb_bottom_output_6_18;
wire wire_sb_bottom_output_6_19;
wire wire_sb_bottom_output_6_2;
wire wire_sb_bottom_output_6_3;
wire wire_sb_bottom_output_6_4;
wire wire_sb_bottom_output_6_5;
wire wire_sb_bottom_output_6_6;
wire wire_sb_bottom_output_6_7;
wire wire_sb_bottom_output_6_8;
wire wire_sb_bottom_output_6_9;
wire wire_sb_bottom_output_7_0;
wire wire_sb_bottom_output_7_1;
wire wire_sb_bottom_output_7_10;
wire wire_sb_bottom_output_7_11;
wire wire_sb_bottom_output_7_12;
wire wire_sb_bottom_output_7_13;
wire wire_sb_bottom_output_7_14;
wire wire_sb_bottom_output_7_15;
wire wire_sb_bottom_output_7_16;
wire wire_sb_bottom_output_7_17;
wire wire_sb_bottom_output_7_18;
wire wire_sb_bottom_output_7_19;
wire wire_sb_bottom_output_7_2;
wire wire_sb_bottom_output_7_3;
wire wire_sb_bottom_output_7_4;
wire wire_sb_bottom_output_7_5;
wire wire_sb_bottom_output_7_6;
wire wire_sb_bottom_output_7_7;
wire wire_sb_bottom_output_7_8;
wire wire_sb_bottom_output_7_9;
wire wire_sb_bottom_output_8_0;
wire wire_sb_bottom_output_8_1;
wire wire_sb_bottom_output_8_10;
wire wire_sb_bottom_output_8_11;
wire wire_sb_bottom_output_8_12;
wire wire_sb_bottom_output_8_13;
wire wire_sb_bottom_output_8_14;
wire wire_sb_bottom_output_8_15;
wire wire_sb_bottom_output_8_16;
wire wire_sb_bottom_output_8_17;
wire wire_sb_bottom_output_8_18;
wire wire_sb_bottom_output_8_19;
wire wire_sb_bottom_output_8_2;
wire wire_sb_bottom_output_8_3;
wire wire_sb_bottom_output_8_4;
wire wire_sb_bottom_output_8_5;
wire wire_sb_bottom_output_8_6;
wire wire_sb_bottom_output_8_7;
wire wire_sb_bottom_output_8_8;
wire wire_sb_bottom_output_8_9;
wire wire_sb_bottom_output_9_0;
wire wire_sb_bottom_output_9_1;
wire wire_sb_bottom_output_9_10;
wire wire_sb_bottom_output_9_11;
wire wire_sb_bottom_output_9_12;
wire wire_sb_bottom_output_9_13;
wire wire_sb_bottom_output_9_14;
wire wire_sb_bottom_output_9_15;
wire wire_sb_bottom_output_9_16;
wire wire_sb_bottom_output_9_17;
wire wire_sb_bottom_output_9_18;
wire wire_sb_bottom_output_9_19;
wire wire_sb_bottom_output_9_2;
wire wire_sb_bottom_output_9_3;
wire wire_sb_bottom_output_9_4;
wire wire_sb_bottom_output_9_5;
wire wire_sb_bottom_output_9_6;
wire wire_sb_bottom_output_9_7;
wire wire_sb_bottom_output_9_8;
wire wire_sb_bottom_output_9_9;
wire wire_sb_left_input_0_0;
wire wire_sb_left_input_0_1;
wire wire_sb_left_input_0_10;
wire wire_sb_left_input_0_11;
wire wire_sb_left_input_0_12;
wire wire_sb_left_input_0_13;
wire wire_sb_left_input_0_14;
wire wire_sb_left_input_0_15;
wire wire_sb_left_input_0_16;
wire wire_sb_left_input_0_17;
wire wire_sb_left_input_0_18;
wire wire_sb_left_input_0_19;
wire wire_sb_left_input_0_2;
wire wire_sb_left_input_0_3;
wire wire_sb_left_input_0_4;
wire wire_sb_left_input_0_5;
wire wire_sb_left_input_0_6;
wire wire_sb_left_input_0_7;
wire wire_sb_left_input_0_8;
wire wire_sb_left_input_0_9;
wire wire_sb_left_input_10_0;
wire wire_sb_left_input_10_1;
wire wire_sb_left_input_10_10;
wire wire_sb_left_input_10_11;
wire wire_sb_left_input_10_12;
wire wire_sb_left_input_10_13;
wire wire_sb_left_input_10_14;
wire wire_sb_left_input_10_15;
wire wire_sb_left_input_10_16;
wire wire_sb_left_input_10_17;
wire wire_sb_left_input_10_18;
wire wire_sb_left_input_10_19;
wire wire_sb_left_input_10_2;
wire wire_sb_left_input_10_3;
wire wire_sb_left_input_10_4;
wire wire_sb_left_input_10_5;
wire wire_sb_left_input_10_6;
wire wire_sb_left_input_10_7;
wire wire_sb_left_input_10_8;
wire wire_sb_left_input_10_9;
wire wire_sb_left_input_11_0;
wire wire_sb_left_input_11_1;
wire wire_sb_left_input_11_10;
wire wire_sb_left_input_11_11;
wire wire_sb_left_input_11_12;
wire wire_sb_left_input_11_13;
wire wire_sb_left_input_11_14;
wire wire_sb_left_input_11_15;
wire wire_sb_left_input_11_16;
wire wire_sb_left_input_11_17;
wire wire_sb_left_input_11_18;
wire wire_sb_left_input_11_19;
wire wire_sb_left_input_11_2;
wire wire_sb_left_input_11_3;
wire wire_sb_left_input_11_4;
wire wire_sb_left_input_11_5;
wire wire_sb_left_input_11_6;
wire wire_sb_left_input_11_7;
wire wire_sb_left_input_11_8;
wire wire_sb_left_input_11_9;
wire wire_sb_left_input_1_0;
wire wire_sb_left_input_1_1;
wire wire_sb_left_input_1_10;
wire wire_sb_left_input_1_11;
wire wire_sb_left_input_1_12;
wire wire_sb_left_input_1_13;
wire wire_sb_left_input_1_14;
wire wire_sb_left_input_1_15;
wire wire_sb_left_input_1_16;
wire wire_sb_left_input_1_17;
wire wire_sb_left_input_1_18;
wire wire_sb_left_input_1_19;
wire wire_sb_left_input_1_2;
wire wire_sb_left_input_1_3;
wire wire_sb_left_input_1_4;
wire wire_sb_left_input_1_5;
wire wire_sb_left_input_1_6;
wire wire_sb_left_input_1_7;
wire wire_sb_left_input_1_8;
wire wire_sb_left_input_1_9;
wire wire_sb_left_input_2_0;
wire wire_sb_left_input_2_1;
wire wire_sb_left_input_2_10;
wire wire_sb_left_input_2_11;
wire wire_sb_left_input_2_12;
wire wire_sb_left_input_2_13;
wire wire_sb_left_input_2_14;
wire wire_sb_left_input_2_15;
wire wire_sb_left_input_2_16;
wire wire_sb_left_input_2_17;
wire wire_sb_left_input_2_18;
wire wire_sb_left_input_2_19;
wire wire_sb_left_input_2_2;
wire wire_sb_left_input_2_3;
wire wire_sb_left_input_2_4;
wire wire_sb_left_input_2_5;
wire wire_sb_left_input_2_6;
wire wire_sb_left_input_2_7;
wire wire_sb_left_input_2_8;
wire wire_sb_left_input_2_9;
wire wire_sb_left_input_3_0;
wire wire_sb_left_input_3_1;
wire wire_sb_left_input_3_10;
wire wire_sb_left_input_3_11;
wire wire_sb_left_input_3_12;
wire wire_sb_left_input_3_13;
wire wire_sb_left_input_3_14;
wire wire_sb_left_input_3_15;
wire wire_sb_left_input_3_16;
wire wire_sb_left_input_3_17;
wire wire_sb_left_input_3_18;
wire wire_sb_left_input_3_19;
wire wire_sb_left_input_3_2;
wire wire_sb_left_input_3_3;
wire wire_sb_left_input_3_4;
wire wire_sb_left_input_3_5;
wire wire_sb_left_input_3_6;
wire wire_sb_left_input_3_7;
wire wire_sb_left_input_3_8;
wire wire_sb_left_input_3_9;
wire wire_sb_left_input_4_0;
wire wire_sb_left_input_4_1;
wire wire_sb_left_input_4_10;
wire wire_sb_left_input_4_11;
wire wire_sb_left_input_4_12;
wire wire_sb_left_input_4_13;
wire wire_sb_left_input_4_14;
wire wire_sb_left_input_4_15;
wire wire_sb_left_input_4_16;
wire wire_sb_left_input_4_17;
wire wire_sb_left_input_4_18;
wire wire_sb_left_input_4_19;
wire wire_sb_left_input_4_2;
wire wire_sb_left_input_4_3;
wire wire_sb_left_input_4_4;
wire wire_sb_left_input_4_5;
wire wire_sb_left_input_4_6;
wire wire_sb_left_input_4_7;
wire wire_sb_left_input_4_8;
wire wire_sb_left_input_4_9;
wire wire_sb_left_input_5_0;
wire wire_sb_left_input_5_1;
wire wire_sb_left_input_5_10;
wire wire_sb_left_input_5_11;
wire wire_sb_left_input_5_12;
wire wire_sb_left_input_5_13;
wire wire_sb_left_input_5_14;
wire wire_sb_left_input_5_15;
wire wire_sb_left_input_5_16;
wire wire_sb_left_input_5_17;
wire wire_sb_left_input_5_18;
wire wire_sb_left_input_5_19;
wire wire_sb_left_input_5_2;
wire wire_sb_left_input_5_3;
wire wire_sb_left_input_5_4;
wire wire_sb_left_input_5_5;
wire wire_sb_left_input_5_6;
wire wire_sb_left_input_5_7;
wire wire_sb_left_input_5_8;
wire wire_sb_left_input_5_9;
wire wire_sb_left_input_6_0;
wire wire_sb_left_input_6_1;
wire wire_sb_left_input_6_10;
wire wire_sb_left_input_6_11;
wire wire_sb_left_input_6_12;
wire wire_sb_left_input_6_13;
wire wire_sb_left_input_6_14;
wire wire_sb_left_input_6_15;
wire wire_sb_left_input_6_16;
wire wire_sb_left_input_6_17;
wire wire_sb_left_input_6_18;
wire wire_sb_left_input_6_19;
wire wire_sb_left_input_6_2;
wire wire_sb_left_input_6_3;
wire wire_sb_left_input_6_4;
wire wire_sb_left_input_6_5;
wire wire_sb_left_input_6_6;
wire wire_sb_left_input_6_7;
wire wire_sb_left_input_6_8;
wire wire_sb_left_input_6_9;
wire wire_sb_left_input_7_0;
wire wire_sb_left_input_7_1;
wire wire_sb_left_input_7_10;
wire wire_sb_left_input_7_11;
wire wire_sb_left_input_7_12;
wire wire_sb_left_input_7_13;
wire wire_sb_left_input_7_14;
wire wire_sb_left_input_7_15;
wire wire_sb_left_input_7_16;
wire wire_sb_left_input_7_17;
wire wire_sb_left_input_7_18;
wire wire_sb_left_input_7_19;
wire wire_sb_left_input_7_2;
wire wire_sb_left_input_7_3;
wire wire_sb_left_input_7_4;
wire wire_sb_left_input_7_5;
wire wire_sb_left_input_7_6;
wire wire_sb_left_input_7_7;
wire wire_sb_left_input_7_8;
wire wire_sb_left_input_7_9;
wire wire_sb_left_input_8_0;
wire wire_sb_left_input_8_1;
wire wire_sb_left_input_8_10;
wire wire_sb_left_input_8_11;
wire wire_sb_left_input_8_12;
wire wire_sb_left_input_8_13;
wire wire_sb_left_input_8_14;
wire wire_sb_left_input_8_15;
wire wire_sb_left_input_8_16;
wire wire_sb_left_input_8_17;
wire wire_sb_left_input_8_18;
wire wire_sb_left_input_8_19;
wire wire_sb_left_input_8_2;
wire wire_sb_left_input_8_3;
wire wire_sb_left_input_8_4;
wire wire_sb_left_input_8_5;
wire wire_sb_left_input_8_6;
wire wire_sb_left_input_8_7;
wire wire_sb_left_input_8_8;
wire wire_sb_left_input_8_9;
wire wire_sb_left_input_9_0;
wire wire_sb_left_input_9_1;
wire wire_sb_left_input_9_10;
wire wire_sb_left_input_9_11;
wire wire_sb_left_input_9_12;
wire wire_sb_left_input_9_13;
wire wire_sb_left_input_9_14;
wire wire_sb_left_input_9_15;
wire wire_sb_left_input_9_16;
wire wire_sb_left_input_9_17;
wire wire_sb_left_input_9_18;
wire wire_sb_left_input_9_19;
wire wire_sb_left_input_9_2;
wire wire_sb_left_input_9_3;
wire wire_sb_left_input_9_4;
wire wire_sb_left_input_9_5;
wire wire_sb_left_input_9_6;
wire wire_sb_left_input_9_7;
wire wire_sb_left_input_9_8;
wire wire_sb_left_input_9_9;
wire wire_sb_left_output_0_0;
wire wire_sb_left_output_0_1;
wire wire_sb_left_output_0_10;
wire wire_sb_left_output_0_11;
wire wire_sb_left_output_0_12;
wire wire_sb_left_output_0_13;
wire wire_sb_left_output_0_14;
wire wire_sb_left_output_0_15;
wire wire_sb_left_output_0_16;
wire wire_sb_left_output_0_17;
wire wire_sb_left_output_0_18;
wire wire_sb_left_output_0_19;
wire wire_sb_left_output_0_2;
wire wire_sb_left_output_0_3;
wire wire_sb_left_output_0_4;
wire wire_sb_left_output_0_5;
wire wire_sb_left_output_0_6;
wire wire_sb_left_output_0_7;
wire wire_sb_left_output_0_8;
wire wire_sb_left_output_0_9;
wire wire_sb_left_output_10_0;
wire wire_sb_left_output_10_1;
wire wire_sb_left_output_10_10;
wire wire_sb_left_output_10_11;
wire wire_sb_left_output_10_12;
wire wire_sb_left_output_10_13;
wire wire_sb_left_output_10_14;
wire wire_sb_left_output_10_15;
wire wire_sb_left_output_10_16;
wire wire_sb_left_output_10_17;
wire wire_sb_left_output_10_18;
wire wire_sb_left_output_10_19;
wire wire_sb_left_output_10_2;
wire wire_sb_left_output_10_3;
wire wire_sb_left_output_10_4;
wire wire_sb_left_output_10_5;
wire wire_sb_left_output_10_6;
wire wire_sb_left_output_10_7;
wire wire_sb_left_output_10_8;
wire wire_sb_left_output_10_9;
wire wire_sb_left_output_11_0;
wire wire_sb_left_output_11_1;
wire wire_sb_left_output_11_10;
wire wire_sb_left_output_11_11;
wire wire_sb_left_output_11_12;
wire wire_sb_left_output_11_13;
wire wire_sb_left_output_11_14;
wire wire_sb_left_output_11_15;
wire wire_sb_left_output_11_16;
wire wire_sb_left_output_11_17;
wire wire_sb_left_output_11_18;
wire wire_sb_left_output_11_19;
wire wire_sb_left_output_11_2;
wire wire_sb_left_output_11_3;
wire wire_sb_left_output_11_4;
wire wire_sb_left_output_11_5;
wire wire_sb_left_output_11_6;
wire wire_sb_left_output_11_7;
wire wire_sb_left_output_11_8;
wire wire_sb_left_output_11_9;
wire wire_sb_left_output_1_0;
wire wire_sb_left_output_1_1;
wire wire_sb_left_output_1_10;
wire wire_sb_left_output_1_11;
wire wire_sb_left_output_1_12;
wire wire_sb_left_output_1_13;
wire wire_sb_left_output_1_14;
wire wire_sb_left_output_1_15;
wire wire_sb_left_output_1_16;
wire wire_sb_left_output_1_17;
wire wire_sb_left_output_1_18;
wire wire_sb_left_output_1_19;
wire wire_sb_left_output_1_2;
wire wire_sb_left_output_1_3;
wire wire_sb_left_output_1_4;
wire wire_sb_left_output_1_5;
wire wire_sb_left_output_1_6;
wire wire_sb_left_output_1_7;
wire wire_sb_left_output_1_8;
wire wire_sb_left_output_1_9;
wire wire_sb_left_output_2_0;
wire wire_sb_left_output_2_1;
wire wire_sb_left_output_2_10;
wire wire_sb_left_output_2_11;
wire wire_sb_left_output_2_12;
wire wire_sb_left_output_2_13;
wire wire_sb_left_output_2_14;
wire wire_sb_left_output_2_15;
wire wire_sb_left_output_2_16;
wire wire_sb_left_output_2_17;
wire wire_sb_left_output_2_18;
wire wire_sb_left_output_2_19;
wire wire_sb_left_output_2_2;
wire wire_sb_left_output_2_3;
wire wire_sb_left_output_2_4;
wire wire_sb_left_output_2_5;
wire wire_sb_left_output_2_6;
wire wire_sb_left_output_2_7;
wire wire_sb_left_output_2_8;
wire wire_sb_left_output_2_9;
wire wire_sb_left_output_3_0;
wire wire_sb_left_output_3_1;
wire wire_sb_left_output_3_10;
wire wire_sb_left_output_3_11;
wire wire_sb_left_output_3_12;
wire wire_sb_left_output_3_13;
wire wire_sb_left_output_3_14;
wire wire_sb_left_output_3_15;
wire wire_sb_left_output_3_16;
wire wire_sb_left_output_3_17;
wire wire_sb_left_output_3_18;
wire wire_sb_left_output_3_19;
wire wire_sb_left_output_3_2;
wire wire_sb_left_output_3_3;
wire wire_sb_left_output_3_4;
wire wire_sb_left_output_3_5;
wire wire_sb_left_output_3_6;
wire wire_sb_left_output_3_7;
wire wire_sb_left_output_3_8;
wire wire_sb_left_output_3_9;
wire wire_sb_left_output_4_0;
wire wire_sb_left_output_4_1;
wire wire_sb_left_output_4_10;
wire wire_sb_left_output_4_11;
wire wire_sb_left_output_4_12;
wire wire_sb_left_output_4_13;
wire wire_sb_left_output_4_14;
wire wire_sb_left_output_4_15;
wire wire_sb_left_output_4_16;
wire wire_sb_left_output_4_17;
wire wire_sb_left_output_4_18;
wire wire_sb_left_output_4_19;
wire wire_sb_left_output_4_2;
wire wire_sb_left_output_4_3;
wire wire_sb_left_output_4_4;
wire wire_sb_left_output_4_5;
wire wire_sb_left_output_4_6;
wire wire_sb_left_output_4_7;
wire wire_sb_left_output_4_8;
wire wire_sb_left_output_4_9;
wire wire_sb_left_output_5_0;
wire wire_sb_left_output_5_1;
wire wire_sb_left_output_5_10;
wire wire_sb_left_output_5_11;
wire wire_sb_left_output_5_12;
wire wire_sb_left_output_5_13;
wire wire_sb_left_output_5_14;
wire wire_sb_left_output_5_15;
wire wire_sb_left_output_5_16;
wire wire_sb_left_output_5_17;
wire wire_sb_left_output_5_18;
wire wire_sb_left_output_5_19;
wire wire_sb_left_output_5_2;
wire wire_sb_left_output_5_3;
wire wire_sb_left_output_5_4;
wire wire_sb_left_output_5_5;
wire wire_sb_left_output_5_6;
wire wire_sb_left_output_5_7;
wire wire_sb_left_output_5_8;
wire wire_sb_left_output_5_9;
wire wire_sb_left_output_6_0;
wire wire_sb_left_output_6_1;
wire wire_sb_left_output_6_10;
wire wire_sb_left_output_6_11;
wire wire_sb_left_output_6_12;
wire wire_sb_left_output_6_13;
wire wire_sb_left_output_6_14;
wire wire_sb_left_output_6_15;
wire wire_sb_left_output_6_16;
wire wire_sb_left_output_6_17;
wire wire_sb_left_output_6_18;
wire wire_sb_left_output_6_19;
wire wire_sb_left_output_6_2;
wire wire_sb_left_output_6_3;
wire wire_sb_left_output_6_4;
wire wire_sb_left_output_6_5;
wire wire_sb_left_output_6_6;
wire wire_sb_left_output_6_7;
wire wire_sb_left_output_6_8;
wire wire_sb_left_output_6_9;
wire wire_sb_left_output_7_0;
wire wire_sb_left_output_7_1;
wire wire_sb_left_output_7_10;
wire wire_sb_left_output_7_11;
wire wire_sb_left_output_7_12;
wire wire_sb_left_output_7_13;
wire wire_sb_left_output_7_14;
wire wire_sb_left_output_7_15;
wire wire_sb_left_output_7_16;
wire wire_sb_left_output_7_17;
wire wire_sb_left_output_7_18;
wire wire_sb_left_output_7_19;
wire wire_sb_left_output_7_2;
wire wire_sb_left_output_7_3;
wire wire_sb_left_output_7_4;
wire wire_sb_left_output_7_5;
wire wire_sb_left_output_7_6;
wire wire_sb_left_output_7_7;
wire wire_sb_left_output_7_8;
wire wire_sb_left_output_7_9;
wire wire_sb_left_output_8_0;
wire wire_sb_left_output_8_1;
wire wire_sb_left_output_8_10;
wire wire_sb_left_output_8_11;
wire wire_sb_left_output_8_12;
wire wire_sb_left_output_8_13;
wire wire_sb_left_output_8_14;
wire wire_sb_left_output_8_15;
wire wire_sb_left_output_8_16;
wire wire_sb_left_output_8_17;
wire wire_sb_left_output_8_18;
wire wire_sb_left_output_8_19;
wire wire_sb_left_output_8_2;
wire wire_sb_left_output_8_3;
wire wire_sb_left_output_8_4;
wire wire_sb_left_output_8_5;
wire wire_sb_left_output_8_6;
wire wire_sb_left_output_8_7;
wire wire_sb_left_output_8_8;
wire wire_sb_left_output_8_9;
wire wire_sb_left_output_9_0;
wire wire_sb_left_output_9_1;
wire wire_sb_left_output_9_10;
wire wire_sb_left_output_9_11;
wire wire_sb_left_output_9_12;
wire wire_sb_left_output_9_13;
wire wire_sb_left_output_9_14;
wire wire_sb_left_output_9_15;
wire wire_sb_left_output_9_16;
wire wire_sb_left_output_9_17;
wire wire_sb_left_output_9_18;
wire wire_sb_left_output_9_19;
wire wire_sb_left_output_9_2;
wire wire_sb_left_output_9_3;
wire wire_sb_left_output_9_4;
wire wire_sb_left_output_9_5;
wire wire_sb_left_output_9_6;
wire wire_sb_left_output_9_7;
wire wire_sb_left_output_9_8;
wire wire_sb_left_output_9_9;
wire [9:0] w_ADDRESS_TILE_0;
wire [24:0] w_SELECT_TILE_0;

loader_mesh_encapsulation loader_mesh_ins(
        .CLK( conf )
      , .RESET( reset )
      , .ADDRESS( { address[14], address[13], address[12], address[11], address[10], address[9], address[8], address[7], address[6], address[5], address[4], address[3], address[2], address[1], address[0] } )
      , .ADDRESS_TILE( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .SELECT_TILE( { w_SELECT_TILE_0[24], w_SELECT_TILE_0[23], w_SELECT_TILE_0[22], w_SELECT_TILE_0[21], w_SELECT_TILE_0[20], w_SELECT_TILE_0[19], w_SELECT_TILE_0[18], w_SELECT_TILE_0[17], w_SELECT_TILE_0[16], w_SELECT_TILE_0[15], w_SELECT_TILE_0[14], w_SELECT_TILE_0[13], w_SELECT_TILE_0[12], w_SELECT_TILE_0[11], w_SELECT_TILE_0[10], w_SELECT_TILE_0[9], w_SELECT_TILE_0[8], w_SELECT_TILE_0[7], w_SELECT_TILE_0[6], w_SELECT_TILE_0[5], w_SELECT_TILE_0[4], w_SELECT_TILE_0[3], w_SELECT_TILE_0[2], w_SELECT_TILE_0[1], w_SELECT_TILE_0[0] } )
     );

TileBoundaryBottom tile_BB21(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[21] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_12, wire_in_cluster_sb_BR_14_12, wire_in_cluster_sb_BR_13_12, wire_in_cluster_sb_BR_12_12, wire_in_cluster_sb_BR_11_12, wire_in_cluster_sb_BR_10_12, wire_in_cluster_sb_BR_9_12, wire_in_cluster_sb_BR_8_12, wire_in_cluster_sb_BR_7_12, wire_in_cluster_sb_BR_6_12, wire_in_cluster_sb_BR_5_12, wire_in_cluster_sb_BR_4_12, wire_in_cluster_sb_BR_3_12, wire_in_cluster_sb_BR_2_12, wire_in_cluster_sb_BR_1_12, wire_in_cluster_sb_BR_0_12 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_13, wire_in_cluster_sb_BL_14_13, wire_in_cluster_sb_BL_13_13, wire_in_cluster_sb_BL_12_13, wire_in_cluster_sb_BL_11_13, wire_in_cluster_sb_BL_10_13, wire_in_cluster_sb_BL_9_13, wire_in_cluster_sb_BL_8_13, wire_in_cluster_sb_BL_7_13, wire_in_cluster_sb_BL_6_13, wire_in_cluster_sb_BL_5_13, wire_in_cluster_sb_BL_4_13, wire_in_cluster_sb_BL_3_13, wire_in_cluster_sb_BL_2_13, wire_in_cluster_sb_BL_1_13, wire_in_cluster_sb_BL_0_13 } )
      , .inpads_0( inpads_bottom[5] )
      , .inpads_1( inpads_bottom[6] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_12, wire_out_cluster_sb_BR_2_12, wire_out_cluster_sb_BR_1_12, wire_out_cluster_sb_BR_0_12 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_13, wire_out_cluster_sb_BL_2_13, wire_out_cluster_sb_BL_1_13, wire_out_cluster_sb_BL_0_13 } )
      , .outpads_0( outpads_bottom[5] )
      , .outpads_1( outpads_bottom[6] )
      , .sb_left_input( { wire_sb_left_input_11_16, wire_sb_left_input_10_16, wire_sb_left_input_9_16, wire_sb_left_input_8_16, wire_sb_left_input_7_16, wire_sb_left_input_6_16, wire_sb_left_input_5_16, wire_sb_left_input_4_16, wire_sb_left_input_3_16, wire_sb_left_input_2_16, wire_sb_left_input_1_16, wire_sb_left_input_0_16 } )
      , .sb_left_output( { wire_sb_left_output_11_16, wire_sb_left_output_10_16, wire_sb_left_output_9_16, wire_sb_left_output_8_16, wire_sb_left_output_7_16, wire_sb_left_output_6_16, wire_sb_left_output_5_16, wire_sb_left_output_4_16, wire_sb_left_output_3_16, wire_sb_left_output_2_16, wire_sb_left_output_1_16, wire_sb_left_output_0_16 } )
      , .sb_right_input( { wire_sb_left_output_11_17, wire_sb_left_output_10_17, wire_sb_left_output_9_17, wire_sb_left_output_8_17, wire_sb_left_output_7_17, wire_sb_left_output_6_17, wire_sb_left_output_5_17, wire_sb_left_output_4_17, wire_sb_left_output_3_17, wire_sb_left_output_2_17, wire_sb_left_output_1_17, wire_sb_left_output_0_17 } )
      , .sb_right_output( { wire_sb_left_input_11_17, wire_sb_left_input_10_17, wire_sb_left_input_9_17, wire_sb_left_input_8_17, wire_sb_left_input_7_17, wire_sb_left_input_6_17, wire_sb_left_input_5_17, wire_sb_left_input_4_17, wire_sb_left_input_3_17, wire_sb_left_input_2_17, wire_sb_left_input_1_17, wire_sb_left_input_0_17 } )
      , .sb_top_input( { wire_sb_bottom_output_11_16, wire_sb_bottom_output_10_16, wire_sb_bottom_output_9_16, wire_sb_bottom_output_8_16, wire_sb_bottom_output_7_16, wire_sb_bottom_output_6_16, wire_sb_bottom_output_5_16, wire_sb_bottom_output_4_16, wire_sb_bottom_output_3_16, wire_sb_bottom_output_2_16, wire_sb_bottom_output_1_16, wire_sb_bottom_output_0_16 } )
      , .sb_top_output( { wire_sb_bottom_input_11_16, wire_sb_bottom_input_10_16, wire_sb_bottom_input_9_16, wire_sb_bottom_input_8_16, wire_sb_bottom_input_7_16, wire_sb_bottom_input_6_16, wire_sb_bottom_input_5_16, wire_sb_bottom_input_4_16, wire_sb_bottom_input_3_16, wire_sb_bottom_input_2_16, wire_sb_bottom_input_1_16, wire_sb_bottom_input_0_16 } )
     );

TileBoundaryBottom tile_BB22(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[22] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_13, wire_in_cluster_sb_BR_14_13, wire_in_cluster_sb_BR_13_13, wire_in_cluster_sb_BR_12_13, wire_in_cluster_sb_BR_11_13, wire_in_cluster_sb_BR_10_13, wire_in_cluster_sb_BR_9_13, wire_in_cluster_sb_BR_8_13, wire_in_cluster_sb_BR_7_13, wire_in_cluster_sb_BR_6_13, wire_in_cluster_sb_BR_5_13, wire_in_cluster_sb_BR_4_13, wire_in_cluster_sb_BR_3_13, wire_in_cluster_sb_BR_2_13, wire_in_cluster_sb_BR_1_13, wire_in_cluster_sb_BR_0_13 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_14, wire_in_cluster_sb_BL_14_14, wire_in_cluster_sb_BL_13_14, wire_in_cluster_sb_BL_12_14, wire_in_cluster_sb_BL_11_14, wire_in_cluster_sb_BL_10_14, wire_in_cluster_sb_BL_9_14, wire_in_cluster_sb_BL_8_14, wire_in_cluster_sb_BL_7_14, wire_in_cluster_sb_BL_6_14, wire_in_cluster_sb_BL_5_14, wire_in_cluster_sb_BL_4_14, wire_in_cluster_sb_BL_3_14, wire_in_cluster_sb_BL_2_14, wire_in_cluster_sb_BL_1_14, wire_in_cluster_sb_BL_0_14 } )
      , .inpads_0( inpads_bottom[3] )
      , .inpads_1( inpads_bottom[4] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_13, wire_out_cluster_sb_BR_2_13, wire_out_cluster_sb_BR_1_13, wire_out_cluster_sb_BR_0_13 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_14, wire_out_cluster_sb_BL_2_14, wire_out_cluster_sb_BL_1_14, wire_out_cluster_sb_BL_0_14 } )
      , .outpads_0( outpads_bottom[3] )
      , .outpads_1( outpads_bottom[4] )
      , .sb_left_input( { wire_sb_left_input_11_17, wire_sb_left_input_10_17, wire_sb_left_input_9_17, wire_sb_left_input_8_17, wire_sb_left_input_7_17, wire_sb_left_input_6_17, wire_sb_left_input_5_17, wire_sb_left_input_4_17, wire_sb_left_input_3_17, wire_sb_left_input_2_17, wire_sb_left_input_1_17, wire_sb_left_input_0_17 } )
      , .sb_left_output( { wire_sb_left_output_11_17, wire_sb_left_output_10_17, wire_sb_left_output_9_17, wire_sb_left_output_8_17, wire_sb_left_output_7_17, wire_sb_left_output_6_17, wire_sb_left_output_5_17, wire_sb_left_output_4_17, wire_sb_left_output_3_17, wire_sb_left_output_2_17, wire_sb_left_output_1_17, wire_sb_left_output_0_17 } )
      , .sb_right_input( { wire_sb_left_output_11_18, wire_sb_left_output_10_18, wire_sb_left_output_9_18, wire_sb_left_output_8_18, wire_sb_left_output_7_18, wire_sb_left_output_6_18, wire_sb_left_output_5_18, wire_sb_left_output_4_18, wire_sb_left_output_3_18, wire_sb_left_output_2_18, wire_sb_left_output_1_18, wire_sb_left_output_0_18 } )
      , .sb_right_output( { wire_sb_left_input_11_18, wire_sb_left_input_10_18, wire_sb_left_input_9_18, wire_sb_left_input_8_18, wire_sb_left_input_7_18, wire_sb_left_input_6_18, wire_sb_left_input_5_18, wire_sb_left_input_4_18, wire_sb_left_input_3_18, wire_sb_left_input_2_18, wire_sb_left_input_1_18, wire_sb_left_input_0_18 } )
      , .sb_top_input( { wire_sb_bottom_output_11_17, wire_sb_bottom_output_10_17, wire_sb_bottom_output_9_17, wire_sb_bottom_output_8_17, wire_sb_bottom_output_7_17, wire_sb_bottom_output_6_17, wire_sb_bottom_output_5_17, wire_sb_bottom_output_4_17, wire_sb_bottom_output_3_17, wire_sb_bottom_output_2_17, wire_sb_bottom_output_1_17, wire_sb_bottom_output_0_17 } )
      , .sb_top_output( { wire_sb_bottom_input_11_17, wire_sb_bottom_input_10_17, wire_sb_bottom_input_9_17, wire_sb_bottom_input_8_17, wire_sb_bottom_input_7_17, wire_sb_bottom_input_6_17, wire_sb_bottom_input_5_17, wire_sb_bottom_input_4_17, wire_sb_bottom_input_3_17, wire_sb_bottom_input_2_17, wire_sb_bottom_input_1_17, wire_sb_bottom_input_0_17 } )
     );

TileBoundaryBottom tile_BB23(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[23] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_14, wire_in_cluster_sb_BR_14_14, wire_in_cluster_sb_BR_13_14, wire_in_cluster_sb_BR_12_14, wire_in_cluster_sb_BR_11_14, wire_in_cluster_sb_BR_10_14, wire_in_cluster_sb_BR_9_14, wire_in_cluster_sb_BR_8_14, wire_in_cluster_sb_BR_7_14, wire_in_cluster_sb_BR_6_14, wire_in_cluster_sb_BR_5_14, wire_in_cluster_sb_BR_4_14, wire_in_cluster_sb_BR_3_14, wire_in_cluster_sb_BR_2_14, wire_in_cluster_sb_BR_1_14, wire_in_cluster_sb_BR_0_14 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_15, wire_in_cluster_sb_BL_14_15, wire_in_cluster_sb_BL_13_15, wire_in_cluster_sb_BL_12_15, wire_in_cluster_sb_BL_11_15, wire_in_cluster_sb_BL_10_15, wire_in_cluster_sb_BL_9_15, wire_in_cluster_sb_BL_8_15, wire_in_cluster_sb_BL_7_15, wire_in_cluster_sb_BL_6_15, wire_in_cluster_sb_BL_5_15, wire_in_cluster_sb_BL_4_15, wire_in_cluster_sb_BL_3_15, wire_in_cluster_sb_BL_2_15, wire_in_cluster_sb_BL_1_15, wire_in_cluster_sb_BL_0_15 } )
      , .inpads_0( inpads_bottom[1] )
      , .inpads_1( inpads_bottom[2] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_14, wire_out_cluster_sb_BR_2_14, wire_out_cluster_sb_BR_1_14, wire_out_cluster_sb_BR_0_14 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_15, wire_out_cluster_sb_BL_2_15, wire_out_cluster_sb_BL_1_15, wire_out_cluster_sb_BL_0_15 } )
      , .outpads_0( outpads_bottom[1] )
      , .outpads_1( outpads_bottom[2] )
      , .sb_left_input( { wire_sb_left_input_11_18, wire_sb_left_input_10_18, wire_sb_left_input_9_18, wire_sb_left_input_8_18, wire_sb_left_input_7_18, wire_sb_left_input_6_18, wire_sb_left_input_5_18, wire_sb_left_input_4_18, wire_sb_left_input_3_18, wire_sb_left_input_2_18, wire_sb_left_input_1_18, wire_sb_left_input_0_18 } )
      , .sb_left_output( { wire_sb_left_output_11_18, wire_sb_left_output_10_18, wire_sb_left_output_9_18, wire_sb_left_output_8_18, wire_sb_left_output_7_18, wire_sb_left_output_6_18, wire_sb_left_output_5_18, wire_sb_left_output_4_18, wire_sb_left_output_3_18, wire_sb_left_output_2_18, wire_sb_left_output_1_18, wire_sb_left_output_0_18 } )
      , .sb_right_input( { wire_sb_left_output_11_19, wire_sb_left_output_10_19, wire_sb_left_output_9_19, wire_sb_left_output_8_19, wire_sb_left_output_7_19, wire_sb_left_output_6_19, wire_sb_left_output_5_19, wire_sb_left_output_4_19, wire_sb_left_output_3_19, wire_sb_left_output_2_19, wire_sb_left_output_1_19, wire_sb_left_output_0_19 } )
      , .sb_right_output( { wire_sb_left_input_11_19, wire_sb_left_input_10_19, wire_sb_left_input_9_19, wire_sb_left_input_8_19, wire_sb_left_input_7_19, wire_sb_left_input_6_19, wire_sb_left_input_5_19, wire_sb_left_input_4_19, wire_sb_left_input_3_19, wire_sb_left_input_2_19, wire_sb_left_input_1_19, wire_sb_left_input_0_19 } )
      , .sb_top_input( { wire_sb_bottom_output_11_18, wire_sb_bottom_output_10_18, wire_sb_bottom_output_9_18, wire_sb_bottom_output_8_18, wire_sb_bottom_output_7_18, wire_sb_bottom_output_6_18, wire_sb_bottom_output_5_18, wire_sb_bottom_output_4_18, wire_sb_bottom_output_3_18, wire_sb_bottom_output_2_18, wire_sb_bottom_output_1_18, wire_sb_bottom_output_0_18 } )
      , .sb_top_output( { wire_sb_bottom_input_11_18, wire_sb_bottom_input_10_18, wire_sb_bottom_input_9_18, wire_sb_bottom_input_8_18, wire_sb_bottom_input_7_18, wire_sb_bottom_input_6_18, wire_sb_bottom_input_5_18, wire_sb_bottom_input_4_18, wire_sb_bottom_input_3_18, wire_sb_bottom_input_2_18, wire_sb_bottom_input_1_18, wire_sb_bottom_input_0_18 } )
     );

TileBoundaryLeft tile_BL10(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[10] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_8, wire_in_cluster_sb_TL_14_8, wire_in_cluster_sb_TL_13_8, wire_in_cluster_sb_TL_12_8, wire_in_cluster_sb_TL_11_8, wire_in_cluster_sb_TL_10_8, wire_in_cluster_sb_TL_9_8, wire_in_cluster_sb_TL_8_8, wire_in_cluster_sb_TL_7_8, wire_in_cluster_sb_TL_6_8, wire_in_cluster_sb_TL_5_8, wire_in_cluster_sb_TL_4_8, wire_in_cluster_sb_TL_3_8, wire_in_cluster_sb_TL_2_8, wire_in_cluster_sb_TL_1_8, wire_in_cluster_sb_TL_0_8 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_4, wire_in_cluster_sb_BL_14_4, wire_in_cluster_sb_BL_13_4, wire_in_cluster_sb_BL_12_4, wire_in_cluster_sb_BL_11_4, wire_in_cluster_sb_BL_10_4, wire_in_cluster_sb_BL_9_4, wire_in_cluster_sb_BL_8_4, wire_in_cluster_sb_BL_7_4, wire_in_cluster_sb_BL_6_4, wire_in_cluster_sb_BL_5_4, wire_in_cluster_sb_BL_4_4, wire_in_cluster_sb_BL_3_4, wire_in_cluster_sb_BL_2_4, wire_in_cluster_sb_BL_1_4, wire_in_cluster_sb_BL_0_4 } )
      , .inpads_0( inpads_left[4] )
      , .inpads_1( inpads_left[3] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_8, wire_out_cluster_sb_TL_2_8, wire_out_cluster_sb_TL_1_8, wire_out_cluster_sb_TL_0_8 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_4, wire_out_cluster_sb_BL_2_4, wire_out_cluster_sb_BL_1_4, wire_out_cluster_sb_BL_0_4 } )
      , .outpads_0( outpads_left[4] )
      , .outpads_1( outpads_left[3] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_10, wire_sb_bottom_input_10_10, wire_sb_bottom_input_9_10, wire_sb_bottom_input_8_10, wire_sb_bottom_input_7_10, wire_sb_bottom_input_6_10, wire_sb_bottom_input_5_10, wire_sb_bottom_input_4_10, wire_sb_bottom_input_3_10, wire_sb_bottom_input_2_10, wire_sb_bottom_input_1_10, wire_sb_bottom_input_0_10 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_10, wire_sb_bottom_output_10_10, wire_sb_bottom_output_9_10, wire_sb_bottom_output_8_10, wire_sb_bottom_output_7_10, wire_sb_bottom_output_6_10, wire_sb_bottom_output_5_10, wire_sb_bottom_output_4_10, wire_sb_bottom_output_3_10, wire_sb_bottom_output_2_10, wire_sb_bottom_output_1_10, wire_sb_bottom_output_0_10 } )
      , .sb_right_input( { wire_sb_left_output_11_8, wire_sb_left_output_10_8, wire_sb_left_output_9_8, wire_sb_left_output_8_8, wire_sb_left_output_7_8, wire_sb_left_output_6_8, wire_sb_left_output_5_8, wire_sb_left_output_4_8, wire_sb_left_output_3_8, wire_sb_left_output_2_8, wire_sb_left_output_1_8, wire_sb_left_output_0_8 } )
      , .sb_right_output( { wire_sb_left_input_11_8, wire_sb_left_input_10_8, wire_sb_left_input_9_8, wire_sb_left_input_8_8, wire_sb_left_input_7_8, wire_sb_left_input_6_8, wire_sb_left_input_5_8, wire_sb_left_input_4_8, wire_sb_left_input_3_8, wire_sb_left_input_2_8, wire_sb_left_input_1_8, wire_sb_left_input_0_8 } )
      , .sb_top_input( { wire_sb_bottom_output_11_5, wire_sb_bottom_output_10_5, wire_sb_bottom_output_9_5, wire_sb_bottom_output_8_5, wire_sb_bottom_output_7_5, wire_sb_bottom_output_6_5, wire_sb_bottom_output_5_5, wire_sb_bottom_output_4_5, wire_sb_bottom_output_3_5, wire_sb_bottom_output_2_5, wire_sb_bottom_output_1_5, wire_sb_bottom_output_0_5 } )
      , .sb_top_output( { wire_sb_bottom_input_11_5, wire_sb_bottom_input_10_5, wire_sb_bottom_input_9_5, wire_sb_bottom_input_8_5, wire_sb_bottom_input_7_5, wire_sb_bottom_input_6_5, wire_sb_bottom_input_5_5, wire_sb_bottom_input_4_5, wire_sb_bottom_input_3_5, wire_sb_bottom_input_2_5, wire_sb_bottom_input_1_5, wire_sb_bottom_input_0_5 } )
     );

TileBoundaryLeft tile_BL15(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[15] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_12, wire_in_cluster_sb_TL_14_12, wire_in_cluster_sb_TL_13_12, wire_in_cluster_sb_TL_12_12, wire_in_cluster_sb_TL_11_12, wire_in_cluster_sb_TL_10_12, wire_in_cluster_sb_TL_9_12, wire_in_cluster_sb_TL_8_12, wire_in_cluster_sb_TL_7_12, wire_in_cluster_sb_TL_6_12, wire_in_cluster_sb_TL_5_12, wire_in_cluster_sb_TL_4_12, wire_in_cluster_sb_TL_3_12, wire_in_cluster_sb_TL_2_12, wire_in_cluster_sb_TL_1_12, wire_in_cluster_sb_TL_0_12 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_8, wire_in_cluster_sb_BL_14_8, wire_in_cluster_sb_BL_13_8, wire_in_cluster_sb_BL_12_8, wire_in_cluster_sb_BL_11_8, wire_in_cluster_sb_BL_10_8, wire_in_cluster_sb_BL_9_8, wire_in_cluster_sb_BL_8_8, wire_in_cluster_sb_BL_7_8, wire_in_cluster_sb_BL_6_8, wire_in_cluster_sb_BL_5_8, wire_in_cluster_sb_BL_4_8, wire_in_cluster_sb_BL_3_8, wire_in_cluster_sb_BL_2_8, wire_in_cluster_sb_BL_1_8, wire_in_cluster_sb_BL_0_8 } )
      , .inpads_0( inpads_left[6] )
      , .inpads_1( inpads_left[5] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_12, wire_out_cluster_sb_TL_2_12, wire_out_cluster_sb_TL_1_12, wire_out_cluster_sb_TL_0_12 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_8, wire_out_cluster_sb_BL_2_8, wire_out_cluster_sb_BL_1_8, wire_out_cluster_sb_BL_0_8 } )
      , .outpads_0( outpads_left[6] )
      , .outpads_1( outpads_left[5] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_15, wire_sb_bottom_input_10_15, wire_sb_bottom_input_9_15, wire_sb_bottom_input_8_15, wire_sb_bottom_input_7_15, wire_sb_bottom_input_6_15, wire_sb_bottom_input_5_15, wire_sb_bottom_input_4_15, wire_sb_bottom_input_3_15, wire_sb_bottom_input_2_15, wire_sb_bottom_input_1_15, wire_sb_bottom_input_0_15 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_15, wire_sb_bottom_output_10_15, wire_sb_bottom_output_9_15, wire_sb_bottom_output_8_15, wire_sb_bottom_output_7_15, wire_sb_bottom_output_6_15, wire_sb_bottom_output_5_15, wire_sb_bottom_output_4_15, wire_sb_bottom_output_3_15, wire_sb_bottom_output_2_15, wire_sb_bottom_output_1_15, wire_sb_bottom_output_0_15 } )
      , .sb_right_input( { wire_sb_left_output_11_12, wire_sb_left_output_10_12, wire_sb_left_output_9_12, wire_sb_left_output_8_12, wire_sb_left_output_7_12, wire_sb_left_output_6_12, wire_sb_left_output_5_12, wire_sb_left_output_4_12, wire_sb_left_output_3_12, wire_sb_left_output_2_12, wire_sb_left_output_1_12, wire_sb_left_output_0_12 } )
      , .sb_right_output( { wire_sb_left_input_11_12, wire_sb_left_input_10_12, wire_sb_left_input_9_12, wire_sb_left_input_8_12, wire_sb_left_input_7_12, wire_sb_left_input_6_12, wire_sb_left_input_5_12, wire_sb_left_input_4_12, wire_sb_left_input_3_12, wire_sb_left_input_2_12, wire_sb_left_input_1_12, wire_sb_left_input_0_12 } )
      , .sb_top_input( { wire_sb_bottom_output_11_10, wire_sb_bottom_output_10_10, wire_sb_bottom_output_9_10, wire_sb_bottom_output_8_10, wire_sb_bottom_output_7_10, wire_sb_bottom_output_6_10, wire_sb_bottom_output_5_10, wire_sb_bottom_output_4_10, wire_sb_bottom_output_3_10, wire_sb_bottom_output_2_10, wire_sb_bottom_output_1_10, wire_sb_bottom_output_0_10 } )
      , .sb_top_output( { wire_sb_bottom_input_11_10, wire_sb_bottom_input_10_10, wire_sb_bottom_input_9_10, wire_sb_bottom_input_8_10, wire_sb_bottom_input_7_10, wire_sb_bottom_input_6_10, wire_sb_bottom_input_5_10, wire_sb_bottom_input_4_10, wire_sb_bottom_input_3_10, wire_sb_bottom_input_2_10, wire_sb_bottom_input_1_10, wire_sb_bottom_input_0_10 } )
     );

TileBoundaryLeft tile_BL5(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[5] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_4, wire_in_cluster_sb_TL_14_4, wire_in_cluster_sb_TL_13_4, wire_in_cluster_sb_TL_12_4, wire_in_cluster_sb_TL_11_4, wire_in_cluster_sb_TL_10_4, wire_in_cluster_sb_TL_9_4, wire_in_cluster_sb_TL_8_4, wire_in_cluster_sb_TL_7_4, wire_in_cluster_sb_TL_6_4, wire_in_cluster_sb_TL_5_4, wire_in_cluster_sb_TL_4_4, wire_in_cluster_sb_TL_3_4, wire_in_cluster_sb_TL_2_4, wire_in_cluster_sb_TL_1_4, wire_in_cluster_sb_TL_0_4 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_0, wire_in_cluster_sb_BL_14_0, wire_in_cluster_sb_BL_13_0, wire_in_cluster_sb_BL_12_0, wire_in_cluster_sb_BL_11_0, wire_in_cluster_sb_BL_10_0, wire_in_cluster_sb_BL_9_0, wire_in_cluster_sb_BL_8_0, wire_in_cluster_sb_BL_7_0, wire_in_cluster_sb_BL_6_0, wire_in_cluster_sb_BL_5_0, wire_in_cluster_sb_BL_4_0, wire_in_cluster_sb_BL_3_0, wire_in_cluster_sb_BL_2_0, wire_in_cluster_sb_BL_1_0, wire_in_cluster_sb_BL_0_0 } )
      , .inpads_0( inpads_left[2] )
      , .inpads_1( inpads_left[1] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_4, wire_out_cluster_sb_TL_2_4, wire_out_cluster_sb_TL_1_4, wire_out_cluster_sb_TL_0_4 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_0, wire_out_cluster_sb_BL_2_0, wire_out_cluster_sb_BL_1_0, wire_out_cluster_sb_BL_0_0 } )
      , .outpads_0( outpads_left[2] )
      , .outpads_1( outpads_left[1] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_5, wire_sb_bottom_input_10_5, wire_sb_bottom_input_9_5, wire_sb_bottom_input_8_5, wire_sb_bottom_input_7_5, wire_sb_bottom_input_6_5, wire_sb_bottom_input_5_5, wire_sb_bottom_input_4_5, wire_sb_bottom_input_3_5, wire_sb_bottom_input_2_5, wire_sb_bottom_input_1_5, wire_sb_bottom_input_0_5 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_5, wire_sb_bottom_output_10_5, wire_sb_bottom_output_9_5, wire_sb_bottom_output_8_5, wire_sb_bottom_output_7_5, wire_sb_bottom_output_6_5, wire_sb_bottom_output_5_5, wire_sb_bottom_output_4_5, wire_sb_bottom_output_3_5, wire_sb_bottom_output_2_5, wire_sb_bottom_output_1_5, wire_sb_bottom_output_0_5 } )
      , .sb_right_input( { wire_sb_left_output_11_4, wire_sb_left_output_10_4, wire_sb_left_output_9_4, wire_sb_left_output_8_4, wire_sb_left_output_7_4, wire_sb_left_output_6_4, wire_sb_left_output_5_4, wire_sb_left_output_4_4, wire_sb_left_output_3_4, wire_sb_left_output_2_4, wire_sb_left_output_1_4, wire_sb_left_output_0_4 } )
      , .sb_right_output( { wire_sb_left_input_11_4, wire_sb_left_input_10_4, wire_sb_left_input_9_4, wire_sb_left_input_8_4, wire_sb_left_input_7_4, wire_sb_left_input_6_4, wire_sb_left_input_5_4, wire_sb_left_input_4_4, wire_sb_left_input_3_4, wire_sb_left_input_2_4, wire_sb_left_input_1_4, wire_sb_left_input_0_4 } )
      , .sb_top_input( { wire_sb_bottom_output_11_0, wire_sb_bottom_output_10_0, wire_sb_bottom_output_9_0, wire_sb_bottom_output_8_0, wire_sb_bottom_output_7_0, wire_sb_bottom_output_6_0, wire_sb_bottom_output_5_0, wire_sb_bottom_output_4_0, wire_sb_bottom_output_3_0, wire_sb_bottom_output_2_0, wire_sb_bottom_output_1_0, wire_sb_bottom_output_0_0 } )
      , .sb_top_output( { wire_sb_bottom_input_11_0, wire_sb_bottom_input_10_0, wire_sb_bottom_input_9_0, wire_sb_bottom_input_8_0, wire_sb_bottom_input_7_0, wire_sb_bottom_input_6_0, wire_sb_bottom_input_5_0, wire_sb_bottom_input_4_0, wire_sb_bottom_input_3_0, wire_sb_bottom_input_2_0, wire_sb_bottom_input_1_0, wire_sb_bottom_input_0_0 } )
     );

TileBoundaryRight tile_BR14(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[14] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_7, wire_in_cluster_sb_BR_14_7, wire_in_cluster_sb_BR_13_7, wire_in_cluster_sb_BR_12_7, wire_in_cluster_sb_BR_11_7, wire_in_cluster_sb_BR_10_7, wire_in_cluster_sb_BR_9_7, wire_in_cluster_sb_BR_8_7, wire_in_cluster_sb_BR_7_7, wire_in_cluster_sb_BR_6_7, wire_in_cluster_sb_BR_5_7, wire_in_cluster_sb_BR_4_7, wire_in_cluster_sb_BR_3_7, wire_in_cluster_sb_BR_2_7, wire_in_cluster_sb_BR_1_7, wire_in_cluster_sb_BR_0_7 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_11, wire_in_cluster_sb_BL_14_11, wire_in_cluster_sb_BL_13_11, wire_in_cluster_sb_BL_12_11, wire_in_cluster_sb_BL_11_11, wire_in_cluster_sb_BL_10_11, wire_in_cluster_sb_BL_9_11, wire_in_cluster_sb_BL_8_11, wire_in_cluster_sb_BL_7_11, wire_in_cluster_sb_BL_6_11, wire_in_cluster_sb_BL_5_11, wire_in_cluster_sb_BL_4_11, wire_in_cluster_sb_BL_3_11, wire_in_cluster_sb_BL_2_11, wire_in_cluster_sb_BL_1_11, wire_in_cluster_sb_BL_0_11 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_11, wire_in_cluster_sb_BR_14_11, wire_in_cluster_sb_BR_13_11, wire_in_cluster_sb_BR_12_11, wire_in_cluster_sb_BR_11_11, wire_in_cluster_sb_BR_10_11, wire_in_cluster_sb_BR_9_11, wire_in_cluster_sb_BR_8_11, wire_in_cluster_sb_BR_7_11, wire_in_cluster_sb_BR_6_11, wire_in_cluster_sb_BR_5_11, wire_in_cluster_sb_BR_4_11, wire_in_cluster_sb_BR_3_11, wire_in_cluster_sb_BR_2_11, wire_in_cluster_sb_BR_1_11, wire_in_cluster_sb_BR_0_11 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_11, wire_in_cluster_sb_TL_14_11, wire_in_cluster_sb_TL_13_11, wire_in_cluster_sb_TL_12_11, wire_in_cluster_sb_TL_11_11, wire_in_cluster_sb_TL_10_11, wire_in_cluster_sb_TL_9_11, wire_in_cluster_sb_TL_8_11, wire_in_cluster_sb_TL_7_11, wire_in_cluster_sb_TL_6_11, wire_in_cluster_sb_TL_5_11, wire_in_cluster_sb_TL_4_11, wire_in_cluster_sb_TL_3_11, wire_in_cluster_sb_TL_2_11, wire_in_cluster_sb_TL_1_11, wire_in_cluster_sb_TL_0_11 } )
      , .inpads_0( inpads_right[3] )
      , .inpads_1( inpads_right[4] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_7, wire_out_cluster_sb_BR_2_7, wire_out_cluster_sb_BR_1_7, wire_out_cluster_sb_BR_0_7 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_11, wire_out_cluster_sb_BL_2_11, wire_out_cluster_sb_BL_1_11, wire_out_cluster_sb_BL_0_11 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_11, wire_out_cluster_sb_BR_2_11, wire_out_cluster_sb_BR_1_11, wire_out_cluster_sb_BR_0_11 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_11, wire_out_cluster_sb_TL_2_11, wire_out_cluster_sb_TL_1_11, wire_out_cluster_sb_TL_0_11 } )
      , .outpads_0( outpads_right[3] )
      , .outpads_1( outpads_right[4] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_14, wire_sb_bottom_input_10_14, wire_sb_bottom_input_9_14, wire_sb_bottom_input_8_14, wire_sb_bottom_input_7_14, wire_sb_bottom_input_6_14, wire_sb_bottom_input_5_14, wire_sb_bottom_input_4_14, wire_sb_bottom_input_3_14, wire_sb_bottom_input_2_14, wire_sb_bottom_input_1_14, wire_sb_bottom_input_0_14 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_14, wire_sb_bottom_output_10_14, wire_sb_bottom_output_9_14, wire_sb_bottom_output_8_14, wire_sb_bottom_output_7_14, wire_sb_bottom_output_6_14, wire_sb_bottom_output_5_14, wire_sb_bottom_output_4_14, wire_sb_bottom_output_3_14, wire_sb_bottom_output_2_14, wire_sb_bottom_output_1_14, wire_sb_bottom_output_0_14 } )
      , .sb_left_input( { wire_sb_left_input_11_11, wire_sb_left_input_10_11, wire_sb_left_input_9_11, wire_sb_left_input_8_11, wire_sb_left_input_7_11, wire_sb_left_input_6_11, wire_sb_left_input_5_11, wire_sb_left_input_4_11, wire_sb_left_input_3_11, wire_sb_left_input_2_11, wire_sb_left_input_1_11, wire_sb_left_input_0_11 } )
      , .sb_left_output( { wire_sb_left_output_11_11, wire_sb_left_output_10_11, wire_sb_left_output_9_11, wire_sb_left_output_8_11, wire_sb_left_output_7_11, wire_sb_left_output_6_11, wire_sb_left_output_5_11, wire_sb_left_output_4_11, wire_sb_left_output_3_11, wire_sb_left_output_2_11, wire_sb_left_output_1_11, wire_sb_left_output_0_11 } )
      , .sb_top_input( { wire_sb_bottom_output_11_9, wire_sb_bottom_output_10_9, wire_sb_bottom_output_9_9, wire_sb_bottom_output_8_9, wire_sb_bottom_output_7_9, wire_sb_bottom_output_6_9, wire_sb_bottom_output_5_9, wire_sb_bottom_output_4_9, wire_sb_bottom_output_3_9, wire_sb_bottom_output_2_9, wire_sb_bottom_output_1_9, wire_sb_bottom_output_0_9 } )
      , .sb_top_output( { wire_sb_bottom_input_11_9, wire_sb_bottom_input_10_9, wire_sb_bottom_input_9_9, wire_sb_bottom_input_8_9, wire_sb_bottom_input_7_9, wire_sb_bottom_input_6_9, wire_sb_bottom_input_5_9, wire_sb_bottom_input_4_9, wire_sb_bottom_input_3_9, wire_sb_bottom_input_2_9, wire_sb_bottom_input_1_9, wire_sb_bottom_input_0_9 } )
     );

TileBoundaryRight tile_BR19(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[19] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_11, wire_in_cluster_sb_BR_14_11, wire_in_cluster_sb_BR_13_11, wire_in_cluster_sb_BR_12_11, wire_in_cluster_sb_BR_11_11, wire_in_cluster_sb_BR_10_11, wire_in_cluster_sb_BR_9_11, wire_in_cluster_sb_BR_8_11, wire_in_cluster_sb_BR_7_11, wire_in_cluster_sb_BR_6_11, wire_in_cluster_sb_BR_5_11, wire_in_cluster_sb_BR_4_11, wire_in_cluster_sb_BR_3_11, wire_in_cluster_sb_BR_2_11, wire_in_cluster_sb_BR_1_11, wire_in_cluster_sb_BR_0_11 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_15, wire_in_cluster_sb_BL_14_15, wire_in_cluster_sb_BL_13_15, wire_in_cluster_sb_BL_12_15, wire_in_cluster_sb_BL_11_15, wire_in_cluster_sb_BL_10_15, wire_in_cluster_sb_BL_9_15, wire_in_cluster_sb_BL_8_15, wire_in_cluster_sb_BL_7_15, wire_in_cluster_sb_BL_6_15, wire_in_cluster_sb_BL_5_15, wire_in_cluster_sb_BL_4_15, wire_in_cluster_sb_BL_3_15, wire_in_cluster_sb_BL_2_15, wire_in_cluster_sb_BL_1_15, wire_in_cluster_sb_BL_0_15 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_15, wire_in_cluster_sb_BR_14_15, wire_in_cluster_sb_BR_13_15, wire_in_cluster_sb_BR_12_15, wire_in_cluster_sb_BR_11_15, wire_in_cluster_sb_BR_10_15, wire_in_cluster_sb_BR_9_15, wire_in_cluster_sb_BR_8_15, wire_in_cluster_sb_BR_7_15, wire_in_cluster_sb_BR_6_15, wire_in_cluster_sb_BR_5_15, wire_in_cluster_sb_BR_4_15, wire_in_cluster_sb_BR_3_15, wire_in_cluster_sb_BR_2_15, wire_in_cluster_sb_BR_1_15, wire_in_cluster_sb_BR_0_15 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_15, wire_in_cluster_sb_TL_14_15, wire_in_cluster_sb_TL_13_15, wire_in_cluster_sb_TL_12_15, wire_in_cluster_sb_TL_11_15, wire_in_cluster_sb_TL_10_15, wire_in_cluster_sb_TL_9_15, wire_in_cluster_sb_TL_8_15, wire_in_cluster_sb_TL_7_15, wire_in_cluster_sb_TL_6_15, wire_in_cluster_sb_TL_5_15, wire_in_cluster_sb_TL_4_15, wire_in_cluster_sb_TL_3_15, wire_in_cluster_sb_TL_2_15, wire_in_cluster_sb_TL_1_15, wire_in_cluster_sb_TL_0_15 } )
      , .inpads_0( inpads_right[5] )
      , .inpads_1( inpads_right[6] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_11, wire_out_cluster_sb_BR_2_11, wire_out_cluster_sb_BR_1_11, wire_out_cluster_sb_BR_0_11 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_15, wire_out_cluster_sb_BL_2_15, wire_out_cluster_sb_BL_1_15, wire_out_cluster_sb_BL_0_15 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_15, wire_out_cluster_sb_BR_2_15, wire_out_cluster_sb_BR_1_15, wire_out_cluster_sb_BR_0_15 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_15, wire_out_cluster_sb_TL_2_15, wire_out_cluster_sb_TL_1_15, wire_out_cluster_sb_TL_0_15 } )
      , .outpads_0( outpads_right[5] )
      , .outpads_1( outpads_right[6] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_19, wire_sb_bottom_input_10_19, wire_sb_bottom_input_9_19, wire_sb_bottom_input_8_19, wire_sb_bottom_input_7_19, wire_sb_bottom_input_6_19, wire_sb_bottom_input_5_19, wire_sb_bottom_input_4_19, wire_sb_bottom_input_3_19, wire_sb_bottom_input_2_19, wire_sb_bottom_input_1_19, wire_sb_bottom_input_0_19 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_19, wire_sb_bottom_output_10_19, wire_sb_bottom_output_9_19, wire_sb_bottom_output_8_19, wire_sb_bottom_output_7_19, wire_sb_bottom_output_6_19, wire_sb_bottom_output_5_19, wire_sb_bottom_output_4_19, wire_sb_bottom_output_3_19, wire_sb_bottom_output_2_19, wire_sb_bottom_output_1_19, wire_sb_bottom_output_0_19 } )
      , .sb_left_input( { wire_sb_left_input_11_15, wire_sb_left_input_10_15, wire_sb_left_input_9_15, wire_sb_left_input_8_15, wire_sb_left_input_7_15, wire_sb_left_input_6_15, wire_sb_left_input_5_15, wire_sb_left_input_4_15, wire_sb_left_input_3_15, wire_sb_left_input_2_15, wire_sb_left_input_1_15, wire_sb_left_input_0_15 } )
      , .sb_left_output( { wire_sb_left_output_11_15, wire_sb_left_output_10_15, wire_sb_left_output_9_15, wire_sb_left_output_8_15, wire_sb_left_output_7_15, wire_sb_left_output_6_15, wire_sb_left_output_5_15, wire_sb_left_output_4_15, wire_sb_left_output_3_15, wire_sb_left_output_2_15, wire_sb_left_output_1_15, wire_sb_left_output_0_15 } )
      , .sb_top_input( { wire_sb_bottom_output_11_14, wire_sb_bottom_output_10_14, wire_sb_bottom_output_9_14, wire_sb_bottom_output_8_14, wire_sb_bottom_output_7_14, wire_sb_bottom_output_6_14, wire_sb_bottom_output_5_14, wire_sb_bottom_output_4_14, wire_sb_bottom_output_3_14, wire_sb_bottom_output_2_14, wire_sb_bottom_output_1_14, wire_sb_bottom_output_0_14 } )
      , .sb_top_output( { wire_sb_bottom_input_11_14, wire_sb_bottom_input_10_14, wire_sb_bottom_input_9_14, wire_sb_bottom_input_8_14, wire_sb_bottom_input_7_14, wire_sb_bottom_input_6_14, wire_sb_bottom_input_5_14, wire_sb_bottom_input_4_14, wire_sb_bottom_input_3_14, wire_sb_bottom_input_2_14, wire_sb_bottom_input_1_14, wire_sb_bottom_input_0_14 } )
     );

TileBoundaryRight tile_BR9(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[9] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_3, wire_in_cluster_sb_BR_14_3, wire_in_cluster_sb_BR_13_3, wire_in_cluster_sb_BR_12_3, wire_in_cluster_sb_BR_11_3, wire_in_cluster_sb_BR_10_3, wire_in_cluster_sb_BR_9_3, wire_in_cluster_sb_BR_8_3, wire_in_cluster_sb_BR_7_3, wire_in_cluster_sb_BR_6_3, wire_in_cluster_sb_BR_5_3, wire_in_cluster_sb_BR_4_3, wire_in_cluster_sb_BR_3_3, wire_in_cluster_sb_BR_2_3, wire_in_cluster_sb_BR_1_3, wire_in_cluster_sb_BR_0_3 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_7, wire_in_cluster_sb_BL_14_7, wire_in_cluster_sb_BL_13_7, wire_in_cluster_sb_BL_12_7, wire_in_cluster_sb_BL_11_7, wire_in_cluster_sb_BL_10_7, wire_in_cluster_sb_BL_9_7, wire_in_cluster_sb_BL_8_7, wire_in_cluster_sb_BL_7_7, wire_in_cluster_sb_BL_6_7, wire_in_cluster_sb_BL_5_7, wire_in_cluster_sb_BL_4_7, wire_in_cluster_sb_BL_3_7, wire_in_cluster_sb_BL_2_7, wire_in_cluster_sb_BL_1_7, wire_in_cluster_sb_BL_0_7 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_7, wire_in_cluster_sb_BR_14_7, wire_in_cluster_sb_BR_13_7, wire_in_cluster_sb_BR_12_7, wire_in_cluster_sb_BR_11_7, wire_in_cluster_sb_BR_10_7, wire_in_cluster_sb_BR_9_7, wire_in_cluster_sb_BR_8_7, wire_in_cluster_sb_BR_7_7, wire_in_cluster_sb_BR_6_7, wire_in_cluster_sb_BR_5_7, wire_in_cluster_sb_BR_4_7, wire_in_cluster_sb_BR_3_7, wire_in_cluster_sb_BR_2_7, wire_in_cluster_sb_BR_1_7, wire_in_cluster_sb_BR_0_7 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_7, wire_in_cluster_sb_TL_14_7, wire_in_cluster_sb_TL_13_7, wire_in_cluster_sb_TL_12_7, wire_in_cluster_sb_TL_11_7, wire_in_cluster_sb_TL_10_7, wire_in_cluster_sb_TL_9_7, wire_in_cluster_sb_TL_8_7, wire_in_cluster_sb_TL_7_7, wire_in_cluster_sb_TL_6_7, wire_in_cluster_sb_TL_5_7, wire_in_cluster_sb_TL_4_7, wire_in_cluster_sb_TL_3_7, wire_in_cluster_sb_TL_2_7, wire_in_cluster_sb_TL_1_7, wire_in_cluster_sb_TL_0_7 } )
      , .inpads_0( inpads_right[1] )
      , .inpads_1( inpads_right[2] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_3, wire_out_cluster_sb_BR_2_3, wire_out_cluster_sb_BR_1_3, wire_out_cluster_sb_BR_0_3 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_7, wire_out_cluster_sb_BL_2_7, wire_out_cluster_sb_BL_1_7, wire_out_cluster_sb_BL_0_7 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_7, wire_out_cluster_sb_BR_2_7, wire_out_cluster_sb_BR_1_7, wire_out_cluster_sb_BR_0_7 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_7, wire_out_cluster_sb_TL_2_7, wire_out_cluster_sb_TL_1_7, wire_out_cluster_sb_TL_0_7 } )
      , .outpads_0( outpads_right[1] )
      , .outpads_1( outpads_right[2] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_9, wire_sb_bottom_input_10_9, wire_sb_bottom_input_9_9, wire_sb_bottom_input_8_9, wire_sb_bottom_input_7_9, wire_sb_bottom_input_6_9, wire_sb_bottom_input_5_9, wire_sb_bottom_input_4_9, wire_sb_bottom_input_3_9, wire_sb_bottom_input_2_9, wire_sb_bottom_input_1_9, wire_sb_bottom_input_0_9 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_9, wire_sb_bottom_output_10_9, wire_sb_bottom_output_9_9, wire_sb_bottom_output_8_9, wire_sb_bottom_output_7_9, wire_sb_bottom_output_6_9, wire_sb_bottom_output_5_9, wire_sb_bottom_output_4_9, wire_sb_bottom_output_3_9, wire_sb_bottom_output_2_9, wire_sb_bottom_output_1_9, wire_sb_bottom_output_0_9 } )
      , .sb_left_input( { wire_sb_left_input_11_7, wire_sb_left_input_10_7, wire_sb_left_input_9_7, wire_sb_left_input_8_7, wire_sb_left_input_7_7, wire_sb_left_input_6_7, wire_sb_left_input_5_7, wire_sb_left_input_4_7, wire_sb_left_input_3_7, wire_sb_left_input_2_7, wire_sb_left_input_1_7, wire_sb_left_input_0_7 } )
      , .sb_left_output( { wire_sb_left_output_11_7, wire_sb_left_output_10_7, wire_sb_left_output_9_7, wire_sb_left_output_8_7, wire_sb_left_output_7_7, wire_sb_left_output_6_7, wire_sb_left_output_5_7, wire_sb_left_output_4_7, wire_sb_left_output_3_7, wire_sb_left_output_2_7, wire_sb_left_output_1_7, wire_sb_left_output_0_7 } )
      , .sb_top_input( { wire_sb_bottom_output_11_4, wire_sb_bottom_output_10_4, wire_sb_bottom_output_9_4, wire_sb_bottom_output_8_4, wire_sb_bottom_output_7_4, wire_sb_bottom_output_6_4, wire_sb_bottom_output_5_4, wire_sb_bottom_output_4_4, wire_sb_bottom_output_3_4, wire_sb_bottom_output_2_4, wire_sb_bottom_output_1_4, wire_sb_bottom_output_0_4 } )
      , .sb_top_output( { wire_sb_bottom_input_11_4, wire_sb_bottom_input_10_4, wire_sb_bottom_input_9_4, wire_sb_bottom_input_8_4, wire_sb_bottom_input_7_4, wire_sb_bottom_input_6_4, wire_sb_bottom_input_5_4, wire_sb_bottom_input_4_4, wire_sb_bottom_input_3_4, wire_sb_bottom_input_2_4, wire_sb_bottom_input_1_4, wire_sb_bottom_input_0_4 } )
     );

TileBoundaryTop tile_BT1(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[1] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_1, wire_in_cluster_sb_TL_14_1, wire_in_cluster_sb_TL_13_1, wire_in_cluster_sb_TL_12_1, wire_in_cluster_sb_TL_11_1, wire_in_cluster_sb_TL_10_1, wire_in_cluster_sb_TL_9_1, wire_in_cluster_sb_TL_8_1, wire_in_cluster_sb_TL_7_1, wire_in_cluster_sb_TL_6_1, wire_in_cluster_sb_TL_5_1, wire_in_cluster_sb_TL_4_1, wire_in_cluster_sb_TL_3_1, wire_in_cluster_sb_TL_2_1, wire_in_cluster_sb_TL_1_1, wire_in_cluster_sb_TL_0_1 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_0, wire_in_cluster_sb_BL_14_0, wire_in_cluster_sb_BL_13_0, wire_in_cluster_sb_BL_12_0, wire_in_cluster_sb_BL_11_0, wire_in_cluster_sb_BL_10_0, wire_in_cluster_sb_BL_9_0, wire_in_cluster_sb_BL_8_0, wire_in_cluster_sb_BL_7_0, wire_in_cluster_sb_BL_6_0, wire_in_cluster_sb_BL_5_0, wire_in_cluster_sb_BL_4_0, wire_in_cluster_sb_BL_3_0, wire_in_cluster_sb_BL_2_0, wire_in_cluster_sb_BL_1_0, wire_in_cluster_sb_BL_0_0 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_0, wire_in_cluster_sb_BR_14_0, wire_in_cluster_sb_BR_13_0, wire_in_cluster_sb_BR_12_0, wire_in_cluster_sb_BR_11_0, wire_in_cluster_sb_BR_10_0, wire_in_cluster_sb_BR_9_0, wire_in_cluster_sb_BR_8_0, wire_in_cluster_sb_BR_7_0, wire_in_cluster_sb_BR_6_0, wire_in_cluster_sb_BR_5_0, wire_in_cluster_sb_BR_4_0, wire_in_cluster_sb_BR_3_0, wire_in_cluster_sb_BR_2_0, wire_in_cluster_sb_BR_1_0, wire_in_cluster_sb_BR_0_0 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_0, wire_in_cluster_sb_TL_14_0, wire_in_cluster_sb_TL_13_0, wire_in_cluster_sb_TL_12_0, wire_in_cluster_sb_TL_11_0, wire_in_cluster_sb_TL_10_0, wire_in_cluster_sb_TL_9_0, wire_in_cluster_sb_TL_8_0, wire_in_cluster_sb_TL_7_0, wire_in_cluster_sb_TL_6_0, wire_in_cluster_sb_TL_5_0, wire_in_cluster_sb_TL_4_0, wire_in_cluster_sb_TL_3_0, wire_in_cluster_sb_TL_2_0, wire_in_cluster_sb_TL_1_0, wire_in_cluster_sb_TL_0_0 } )
      , .inpads_0( inpads_top[5] )
      , .inpads_1( inpads_top[6] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_1, wire_out_cluster_sb_TL_2_1, wire_out_cluster_sb_TL_1_1, wire_out_cluster_sb_TL_0_1 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_0, wire_out_cluster_sb_BL_2_0, wire_out_cluster_sb_BL_1_0, wire_out_cluster_sb_BL_0_0 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_0, wire_out_cluster_sb_BR_2_0, wire_out_cluster_sb_BR_1_0, wire_out_cluster_sb_BR_0_0 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_0, wire_out_cluster_sb_TL_2_0, wire_out_cluster_sb_TL_1_0, wire_out_cluster_sb_TL_0_0 } )
      , .outpads_0( outpads_top[5] )
      , .outpads_1( outpads_top[6] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_1, wire_sb_bottom_input_10_1, wire_sb_bottom_input_9_1, wire_sb_bottom_input_8_1, wire_sb_bottom_input_7_1, wire_sb_bottom_input_6_1, wire_sb_bottom_input_5_1, wire_sb_bottom_input_4_1, wire_sb_bottom_input_3_1, wire_sb_bottom_input_2_1, wire_sb_bottom_input_1_1, wire_sb_bottom_input_0_1 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_1, wire_sb_bottom_output_10_1, wire_sb_bottom_output_9_1, wire_sb_bottom_output_8_1, wire_sb_bottom_output_7_1, wire_sb_bottom_output_6_1, wire_sb_bottom_output_5_1, wire_sb_bottom_output_4_1, wire_sb_bottom_output_3_1, wire_sb_bottom_output_2_1, wire_sb_bottom_output_1_1, wire_sb_bottom_output_0_1 } )
      , .sb_left_input( { wire_sb_left_input_11_0, wire_sb_left_input_10_0, wire_sb_left_input_9_0, wire_sb_left_input_8_0, wire_sb_left_input_7_0, wire_sb_left_input_6_0, wire_sb_left_input_5_0, wire_sb_left_input_4_0, wire_sb_left_input_3_0, wire_sb_left_input_2_0, wire_sb_left_input_1_0, wire_sb_left_input_0_0 } )
      , .sb_left_output( { wire_sb_left_output_11_0, wire_sb_left_output_10_0, wire_sb_left_output_9_0, wire_sb_left_output_8_0, wire_sb_left_output_7_0, wire_sb_left_output_6_0, wire_sb_left_output_5_0, wire_sb_left_output_4_0, wire_sb_left_output_3_0, wire_sb_left_output_2_0, wire_sb_left_output_1_0, wire_sb_left_output_0_0 } )
      , .sb_right_input( { wire_sb_left_output_11_1, wire_sb_left_output_10_1, wire_sb_left_output_9_1, wire_sb_left_output_8_1, wire_sb_left_output_7_1, wire_sb_left_output_6_1, wire_sb_left_output_5_1, wire_sb_left_output_4_1, wire_sb_left_output_3_1, wire_sb_left_output_2_1, wire_sb_left_output_1_1, wire_sb_left_output_0_1 } )
      , .sb_right_output( { wire_sb_left_input_11_1, wire_sb_left_input_10_1, wire_sb_left_input_9_1, wire_sb_left_input_8_1, wire_sb_left_input_7_1, wire_sb_left_input_6_1, wire_sb_left_input_5_1, wire_sb_left_input_4_1, wire_sb_left_input_3_1, wire_sb_left_input_2_1, wire_sb_left_input_1_1, wire_sb_left_input_0_1 } )
     );

TileBoundaryTop tile_BT2(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[2] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_2, wire_in_cluster_sb_TL_14_2, wire_in_cluster_sb_TL_13_2, wire_in_cluster_sb_TL_12_2, wire_in_cluster_sb_TL_11_2, wire_in_cluster_sb_TL_10_2, wire_in_cluster_sb_TL_9_2, wire_in_cluster_sb_TL_8_2, wire_in_cluster_sb_TL_7_2, wire_in_cluster_sb_TL_6_2, wire_in_cluster_sb_TL_5_2, wire_in_cluster_sb_TL_4_2, wire_in_cluster_sb_TL_3_2, wire_in_cluster_sb_TL_2_2, wire_in_cluster_sb_TL_1_2, wire_in_cluster_sb_TL_0_2 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_1, wire_in_cluster_sb_BL_14_1, wire_in_cluster_sb_BL_13_1, wire_in_cluster_sb_BL_12_1, wire_in_cluster_sb_BL_11_1, wire_in_cluster_sb_BL_10_1, wire_in_cluster_sb_BL_9_1, wire_in_cluster_sb_BL_8_1, wire_in_cluster_sb_BL_7_1, wire_in_cluster_sb_BL_6_1, wire_in_cluster_sb_BL_5_1, wire_in_cluster_sb_BL_4_1, wire_in_cluster_sb_BL_3_1, wire_in_cluster_sb_BL_2_1, wire_in_cluster_sb_BL_1_1, wire_in_cluster_sb_BL_0_1 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_1, wire_in_cluster_sb_BR_14_1, wire_in_cluster_sb_BR_13_1, wire_in_cluster_sb_BR_12_1, wire_in_cluster_sb_BR_11_1, wire_in_cluster_sb_BR_10_1, wire_in_cluster_sb_BR_9_1, wire_in_cluster_sb_BR_8_1, wire_in_cluster_sb_BR_7_1, wire_in_cluster_sb_BR_6_1, wire_in_cluster_sb_BR_5_1, wire_in_cluster_sb_BR_4_1, wire_in_cluster_sb_BR_3_1, wire_in_cluster_sb_BR_2_1, wire_in_cluster_sb_BR_1_1, wire_in_cluster_sb_BR_0_1 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_1, wire_in_cluster_sb_TL_14_1, wire_in_cluster_sb_TL_13_1, wire_in_cluster_sb_TL_12_1, wire_in_cluster_sb_TL_11_1, wire_in_cluster_sb_TL_10_1, wire_in_cluster_sb_TL_9_1, wire_in_cluster_sb_TL_8_1, wire_in_cluster_sb_TL_7_1, wire_in_cluster_sb_TL_6_1, wire_in_cluster_sb_TL_5_1, wire_in_cluster_sb_TL_4_1, wire_in_cluster_sb_TL_3_1, wire_in_cluster_sb_TL_2_1, wire_in_cluster_sb_TL_1_1, wire_in_cluster_sb_TL_0_1 } )
      , .inpads_0( inpads_top[3] )
      , .inpads_1( inpads_top[4] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_2, wire_out_cluster_sb_TL_2_2, wire_out_cluster_sb_TL_1_2, wire_out_cluster_sb_TL_0_2 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_1, wire_out_cluster_sb_BL_2_1, wire_out_cluster_sb_BL_1_1, wire_out_cluster_sb_BL_0_1 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_1, wire_out_cluster_sb_BR_2_1, wire_out_cluster_sb_BR_1_1, wire_out_cluster_sb_BR_0_1 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_1, wire_out_cluster_sb_TL_2_1, wire_out_cluster_sb_TL_1_1, wire_out_cluster_sb_TL_0_1 } )
      , .outpads_0( outpads_top[3] )
      , .outpads_1( outpads_top[4] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_2, wire_sb_bottom_input_10_2, wire_sb_bottom_input_9_2, wire_sb_bottom_input_8_2, wire_sb_bottom_input_7_2, wire_sb_bottom_input_6_2, wire_sb_bottom_input_5_2, wire_sb_bottom_input_4_2, wire_sb_bottom_input_3_2, wire_sb_bottom_input_2_2, wire_sb_bottom_input_1_2, wire_sb_bottom_input_0_2 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_2, wire_sb_bottom_output_10_2, wire_sb_bottom_output_9_2, wire_sb_bottom_output_8_2, wire_sb_bottom_output_7_2, wire_sb_bottom_output_6_2, wire_sb_bottom_output_5_2, wire_sb_bottom_output_4_2, wire_sb_bottom_output_3_2, wire_sb_bottom_output_2_2, wire_sb_bottom_output_1_2, wire_sb_bottom_output_0_2 } )
      , .sb_left_input( { wire_sb_left_input_11_1, wire_sb_left_input_10_1, wire_sb_left_input_9_1, wire_sb_left_input_8_1, wire_sb_left_input_7_1, wire_sb_left_input_6_1, wire_sb_left_input_5_1, wire_sb_left_input_4_1, wire_sb_left_input_3_1, wire_sb_left_input_2_1, wire_sb_left_input_1_1, wire_sb_left_input_0_1 } )
      , .sb_left_output( { wire_sb_left_output_11_1, wire_sb_left_output_10_1, wire_sb_left_output_9_1, wire_sb_left_output_8_1, wire_sb_left_output_7_1, wire_sb_left_output_6_1, wire_sb_left_output_5_1, wire_sb_left_output_4_1, wire_sb_left_output_3_1, wire_sb_left_output_2_1, wire_sb_left_output_1_1, wire_sb_left_output_0_1 } )
      , .sb_right_input( { wire_sb_left_output_11_2, wire_sb_left_output_10_2, wire_sb_left_output_9_2, wire_sb_left_output_8_2, wire_sb_left_output_7_2, wire_sb_left_output_6_2, wire_sb_left_output_5_2, wire_sb_left_output_4_2, wire_sb_left_output_3_2, wire_sb_left_output_2_2, wire_sb_left_output_1_2, wire_sb_left_output_0_2 } )
      , .sb_right_output( { wire_sb_left_input_11_2, wire_sb_left_input_10_2, wire_sb_left_input_9_2, wire_sb_left_input_8_2, wire_sb_left_input_7_2, wire_sb_left_input_6_2, wire_sb_left_input_5_2, wire_sb_left_input_4_2, wire_sb_left_input_3_2, wire_sb_left_input_2_2, wire_sb_left_input_1_2, wire_sb_left_input_0_2 } )
     );

TileBoundaryTop tile_BT3(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[3] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_3, wire_in_cluster_sb_TL_14_3, wire_in_cluster_sb_TL_13_3, wire_in_cluster_sb_TL_12_3, wire_in_cluster_sb_TL_11_3, wire_in_cluster_sb_TL_10_3, wire_in_cluster_sb_TL_9_3, wire_in_cluster_sb_TL_8_3, wire_in_cluster_sb_TL_7_3, wire_in_cluster_sb_TL_6_3, wire_in_cluster_sb_TL_5_3, wire_in_cluster_sb_TL_4_3, wire_in_cluster_sb_TL_3_3, wire_in_cluster_sb_TL_2_3, wire_in_cluster_sb_TL_1_3, wire_in_cluster_sb_TL_0_3 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_2, wire_in_cluster_sb_BL_14_2, wire_in_cluster_sb_BL_13_2, wire_in_cluster_sb_BL_12_2, wire_in_cluster_sb_BL_11_2, wire_in_cluster_sb_BL_10_2, wire_in_cluster_sb_BL_9_2, wire_in_cluster_sb_BL_8_2, wire_in_cluster_sb_BL_7_2, wire_in_cluster_sb_BL_6_2, wire_in_cluster_sb_BL_5_2, wire_in_cluster_sb_BL_4_2, wire_in_cluster_sb_BL_3_2, wire_in_cluster_sb_BL_2_2, wire_in_cluster_sb_BL_1_2, wire_in_cluster_sb_BL_0_2 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_2, wire_in_cluster_sb_BR_14_2, wire_in_cluster_sb_BR_13_2, wire_in_cluster_sb_BR_12_2, wire_in_cluster_sb_BR_11_2, wire_in_cluster_sb_BR_10_2, wire_in_cluster_sb_BR_9_2, wire_in_cluster_sb_BR_8_2, wire_in_cluster_sb_BR_7_2, wire_in_cluster_sb_BR_6_2, wire_in_cluster_sb_BR_5_2, wire_in_cluster_sb_BR_4_2, wire_in_cluster_sb_BR_3_2, wire_in_cluster_sb_BR_2_2, wire_in_cluster_sb_BR_1_2, wire_in_cluster_sb_BR_0_2 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_2, wire_in_cluster_sb_TL_14_2, wire_in_cluster_sb_TL_13_2, wire_in_cluster_sb_TL_12_2, wire_in_cluster_sb_TL_11_2, wire_in_cluster_sb_TL_10_2, wire_in_cluster_sb_TL_9_2, wire_in_cluster_sb_TL_8_2, wire_in_cluster_sb_TL_7_2, wire_in_cluster_sb_TL_6_2, wire_in_cluster_sb_TL_5_2, wire_in_cluster_sb_TL_4_2, wire_in_cluster_sb_TL_3_2, wire_in_cluster_sb_TL_2_2, wire_in_cluster_sb_TL_1_2, wire_in_cluster_sb_TL_0_2 } )
      , .inpads_0( inpads_top[1] )
      , .inpads_1( inpads_top[2] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_3, wire_out_cluster_sb_TL_2_3, wire_out_cluster_sb_TL_1_3, wire_out_cluster_sb_TL_0_3 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_2, wire_out_cluster_sb_BL_2_2, wire_out_cluster_sb_BL_1_2, wire_out_cluster_sb_BL_0_2 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_2, wire_out_cluster_sb_BR_2_2, wire_out_cluster_sb_BR_1_2, wire_out_cluster_sb_BR_0_2 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_2, wire_out_cluster_sb_TL_2_2, wire_out_cluster_sb_TL_1_2, wire_out_cluster_sb_TL_0_2 } )
      , .outpads_0( outpads_top[1] )
      , .outpads_1( outpads_top[2] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_3, wire_sb_bottom_input_10_3, wire_sb_bottom_input_9_3, wire_sb_bottom_input_8_3, wire_sb_bottom_input_7_3, wire_sb_bottom_input_6_3, wire_sb_bottom_input_5_3, wire_sb_bottom_input_4_3, wire_sb_bottom_input_3_3, wire_sb_bottom_input_2_3, wire_sb_bottom_input_1_3, wire_sb_bottom_input_0_3 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_3, wire_sb_bottom_output_10_3, wire_sb_bottom_output_9_3, wire_sb_bottom_output_8_3, wire_sb_bottom_output_7_3, wire_sb_bottom_output_6_3, wire_sb_bottom_output_5_3, wire_sb_bottom_output_4_3, wire_sb_bottom_output_3_3, wire_sb_bottom_output_2_3, wire_sb_bottom_output_1_3, wire_sb_bottom_output_0_3 } )
      , .sb_left_input( { wire_sb_left_input_11_2, wire_sb_left_input_10_2, wire_sb_left_input_9_2, wire_sb_left_input_8_2, wire_sb_left_input_7_2, wire_sb_left_input_6_2, wire_sb_left_input_5_2, wire_sb_left_input_4_2, wire_sb_left_input_3_2, wire_sb_left_input_2_2, wire_sb_left_input_1_2, wire_sb_left_input_0_2 } )
      , .sb_left_output( { wire_sb_left_output_11_2, wire_sb_left_output_10_2, wire_sb_left_output_9_2, wire_sb_left_output_8_2, wire_sb_left_output_7_2, wire_sb_left_output_6_2, wire_sb_left_output_5_2, wire_sb_left_output_4_2, wire_sb_left_output_3_2, wire_sb_left_output_2_2, wire_sb_left_output_1_2, wire_sb_left_output_0_2 } )
      , .sb_right_input( { wire_sb_left_output_11_3, wire_sb_left_output_10_3, wire_sb_left_output_9_3, wire_sb_left_output_8_3, wire_sb_left_output_7_3, wire_sb_left_output_6_3, wire_sb_left_output_5_3, wire_sb_left_output_4_3, wire_sb_left_output_3_3, wire_sb_left_output_2_3, wire_sb_left_output_1_3, wire_sb_left_output_0_3 } )
      , .sb_right_output( { wire_sb_left_input_11_3, wire_sb_left_input_10_3, wire_sb_left_input_9_3, wire_sb_left_input_8_3, wire_sb_left_input_7_3, wire_sb_left_input_6_3, wire_sb_left_input_5_3, wire_sb_left_input_4_3, wire_sb_left_input_3_3, wire_sb_left_input_2_3, wire_sb_left_input_1_3, wire_sb_left_input_0_3 } )
     );

TileCornerBottomLeft tile_CBL20(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[20] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_12, wire_in_cluster_sb_BL_14_12, wire_in_cluster_sb_BL_13_12, wire_in_cluster_sb_BL_12_12, wire_in_cluster_sb_BL_11_12, wire_in_cluster_sb_BL_10_12, wire_in_cluster_sb_BL_9_12, wire_in_cluster_sb_BL_8_12, wire_in_cluster_sb_BL_7_12, wire_in_cluster_sb_BL_6_12, wire_in_cluster_sb_BL_5_12, wire_in_cluster_sb_BL_4_12, wire_in_cluster_sb_BL_3_12, wire_in_cluster_sb_BL_2_12, wire_in_cluster_sb_BL_1_12, wire_in_cluster_sb_BL_0_12 } )
      , .inpads_0( inpads_bottom[7] )
      , .inpads_1( inpads_left[7] )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_12, wire_out_cluster_sb_BL_2_12, wire_out_cluster_sb_BL_1_12, wire_out_cluster_sb_BL_0_12 } )
      , .outpads_0( outpads_bottom[7] )
      , .outpads_1( outpads_left[7] )
      , .sb_right_input( { wire_sb_left_output_11_16, wire_sb_left_output_10_16, wire_sb_left_output_9_16, wire_sb_left_output_8_16, wire_sb_left_output_7_16, wire_sb_left_output_6_16, wire_sb_left_output_5_16, wire_sb_left_output_4_16, wire_sb_left_output_3_16, wire_sb_left_output_2_16, wire_sb_left_output_1_16, wire_sb_left_output_0_16 } )
      , .sb_right_output( { wire_sb_left_input_11_16, wire_sb_left_input_10_16, wire_sb_left_input_9_16, wire_sb_left_input_8_16, wire_sb_left_input_7_16, wire_sb_left_input_6_16, wire_sb_left_input_5_16, wire_sb_left_input_4_16, wire_sb_left_input_3_16, wire_sb_left_input_2_16, wire_sb_left_input_1_16, wire_sb_left_input_0_16 } )
      , .sb_top_input( { wire_sb_bottom_output_11_15, wire_sb_bottom_output_10_15, wire_sb_bottom_output_9_15, wire_sb_bottom_output_8_15, wire_sb_bottom_output_7_15, wire_sb_bottom_output_6_15, wire_sb_bottom_output_5_15, wire_sb_bottom_output_4_15, wire_sb_bottom_output_3_15, wire_sb_bottom_output_2_15, wire_sb_bottom_output_1_15, wire_sb_bottom_output_0_15 } )
      , .sb_top_output( { wire_sb_bottom_input_11_15, wire_sb_bottom_input_10_15, wire_sb_bottom_input_9_15, wire_sb_bottom_input_8_15, wire_sb_bottom_input_7_15, wire_sb_bottom_input_6_15, wire_sb_bottom_input_5_15, wire_sb_bottom_input_4_15, wire_sb_bottom_input_3_15, wire_sb_bottom_input_2_15, wire_sb_bottom_input_1_15, wire_sb_bottom_input_0_15 } )
     );

TileCornerBottomRight tile_CBR24(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[24] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_15, wire_in_cluster_sb_BR_14_15, wire_in_cluster_sb_BR_13_15, wire_in_cluster_sb_BR_12_15, wire_in_cluster_sb_BR_11_15, wire_in_cluster_sb_BR_10_15, wire_in_cluster_sb_BR_9_15, wire_in_cluster_sb_BR_8_15, wire_in_cluster_sb_BR_7_15, wire_in_cluster_sb_BR_6_15, wire_in_cluster_sb_BR_5_15, wire_in_cluster_sb_BR_4_15, wire_in_cluster_sb_BR_3_15, wire_in_cluster_sb_BR_2_15, wire_in_cluster_sb_BR_1_15, wire_in_cluster_sb_BR_0_15 } )
      , .inpads_0( inpads_right[7] )
      , .inpads_1( inpads_bottom[0] )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_15, wire_out_cluster_sb_BR_2_15, wire_out_cluster_sb_BR_1_15, wire_out_cluster_sb_BR_0_15 } )
      , .outpads_0( outpads_right[7] )
      , .outpads_1( outpads_bottom[0] )
      , .sb_left_input( { wire_sb_left_input_11_19, wire_sb_left_input_10_19, wire_sb_left_input_9_19, wire_sb_left_input_8_19, wire_sb_left_input_7_19, wire_sb_left_input_6_19, wire_sb_left_input_5_19, wire_sb_left_input_4_19, wire_sb_left_input_3_19, wire_sb_left_input_2_19, wire_sb_left_input_1_19, wire_sb_left_input_0_19 } )
      , .sb_left_output( { wire_sb_left_output_11_19, wire_sb_left_output_10_19, wire_sb_left_output_9_19, wire_sb_left_output_8_19, wire_sb_left_output_7_19, wire_sb_left_output_6_19, wire_sb_left_output_5_19, wire_sb_left_output_4_19, wire_sb_left_output_3_19, wire_sb_left_output_2_19, wire_sb_left_output_1_19, wire_sb_left_output_0_19 } )
      , .sb_top_input( { wire_sb_bottom_output_11_19, wire_sb_bottom_output_10_19, wire_sb_bottom_output_9_19, wire_sb_bottom_output_8_19, wire_sb_bottom_output_7_19, wire_sb_bottom_output_6_19, wire_sb_bottom_output_5_19, wire_sb_bottom_output_4_19, wire_sb_bottom_output_3_19, wire_sb_bottom_output_2_19, wire_sb_bottom_output_1_19, wire_sb_bottom_output_0_19 } )
      , .sb_top_output( { wire_sb_bottom_input_11_19, wire_sb_bottom_input_10_19, wire_sb_bottom_input_9_19, wire_sb_bottom_input_8_19, wire_sb_bottom_input_7_19, wire_sb_bottom_input_6_19, wire_sb_bottom_input_5_19, wire_sb_bottom_input_4_19, wire_sb_bottom_input_3_19, wire_sb_bottom_input_2_19, wire_sb_bottom_input_1_19, wire_sb_bottom_input_0_19 } )
     );

TileCornerTopLeft tile_CTL0(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[0] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_0, wire_in_cluster_sb_TL_14_0, wire_in_cluster_sb_TL_13_0, wire_in_cluster_sb_TL_12_0, wire_in_cluster_sb_TL_11_0, wire_in_cluster_sb_TL_10_0, wire_in_cluster_sb_TL_9_0, wire_in_cluster_sb_TL_8_0, wire_in_cluster_sb_TL_7_0, wire_in_cluster_sb_TL_6_0, wire_in_cluster_sb_TL_5_0, wire_in_cluster_sb_TL_4_0, wire_in_cluster_sb_TL_3_0, wire_in_cluster_sb_TL_2_0, wire_in_cluster_sb_TL_1_0, wire_in_cluster_sb_TL_0_0 } )
      , .inpads_0( inpads_top[7] )
      , .inpads_1( inpads_left[0] )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_0, wire_out_cluster_sb_TL_2_0, wire_out_cluster_sb_TL_1_0, wire_out_cluster_sb_TL_0_0 } )
      , .outpads_0( outpads_top[7] )
      , .outpads_1( outpads_left[0] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_0, wire_sb_bottom_input_10_0, wire_sb_bottom_input_9_0, wire_sb_bottom_input_8_0, wire_sb_bottom_input_7_0, wire_sb_bottom_input_6_0, wire_sb_bottom_input_5_0, wire_sb_bottom_input_4_0, wire_sb_bottom_input_3_0, wire_sb_bottom_input_2_0, wire_sb_bottom_input_1_0, wire_sb_bottom_input_0_0 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_0, wire_sb_bottom_output_10_0, wire_sb_bottom_output_9_0, wire_sb_bottom_output_8_0, wire_sb_bottom_output_7_0, wire_sb_bottom_output_6_0, wire_sb_bottom_output_5_0, wire_sb_bottom_output_4_0, wire_sb_bottom_output_3_0, wire_sb_bottom_output_2_0, wire_sb_bottom_output_1_0, wire_sb_bottom_output_0_0 } )
      , .sb_right_input( { wire_sb_left_output_11_0, wire_sb_left_output_10_0, wire_sb_left_output_9_0, wire_sb_left_output_8_0, wire_sb_left_output_7_0, wire_sb_left_output_6_0, wire_sb_left_output_5_0, wire_sb_left_output_4_0, wire_sb_left_output_3_0, wire_sb_left_output_2_0, wire_sb_left_output_1_0, wire_sb_left_output_0_0 } )
      , .sb_right_output( { wire_sb_left_input_11_0, wire_sb_left_input_10_0, wire_sb_left_input_9_0, wire_sb_left_input_8_0, wire_sb_left_input_7_0, wire_sb_left_input_6_0, wire_sb_left_input_5_0, wire_sb_left_input_4_0, wire_sb_left_input_3_0, wire_sb_left_input_2_0, wire_sb_left_input_1_0, wire_sb_left_input_0_0 } )
     );

TileCornerTopRight tile_CTR4(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[4] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_3, wire_in_cluster_sb_BL_14_3, wire_in_cluster_sb_BL_13_3, wire_in_cluster_sb_BL_12_3, wire_in_cluster_sb_BL_11_3, wire_in_cluster_sb_BL_10_3, wire_in_cluster_sb_BL_9_3, wire_in_cluster_sb_BL_8_3, wire_in_cluster_sb_BL_7_3, wire_in_cluster_sb_BL_6_3, wire_in_cluster_sb_BL_5_3, wire_in_cluster_sb_BL_4_3, wire_in_cluster_sb_BL_3_3, wire_in_cluster_sb_BL_2_3, wire_in_cluster_sb_BL_1_3, wire_in_cluster_sb_BL_0_3 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_3, wire_in_cluster_sb_BR_14_3, wire_in_cluster_sb_BR_13_3, wire_in_cluster_sb_BR_12_3, wire_in_cluster_sb_BR_11_3, wire_in_cluster_sb_BR_10_3, wire_in_cluster_sb_BR_9_3, wire_in_cluster_sb_BR_8_3, wire_in_cluster_sb_BR_7_3, wire_in_cluster_sb_BR_6_3, wire_in_cluster_sb_BR_5_3, wire_in_cluster_sb_BR_4_3, wire_in_cluster_sb_BR_3_3, wire_in_cluster_sb_BR_2_3, wire_in_cluster_sb_BR_1_3, wire_in_cluster_sb_BR_0_3 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_3, wire_in_cluster_sb_TL_14_3, wire_in_cluster_sb_TL_13_3, wire_in_cluster_sb_TL_12_3, wire_in_cluster_sb_TL_11_3, wire_in_cluster_sb_TL_10_3, wire_in_cluster_sb_TL_9_3, wire_in_cluster_sb_TL_8_3, wire_in_cluster_sb_TL_7_3, wire_in_cluster_sb_TL_6_3, wire_in_cluster_sb_TL_5_3, wire_in_cluster_sb_TL_4_3, wire_in_cluster_sb_TL_3_3, wire_in_cluster_sb_TL_2_3, wire_in_cluster_sb_TL_1_3, wire_in_cluster_sb_TL_0_3 } )
      , .inpads_0( inpads_right[0] )
      , .inpads_1( inpads_top[0] )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_3, wire_out_cluster_sb_BL_2_3, wire_out_cluster_sb_BL_1_3, wire_out_cluster_sb_BL_0_3 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_3, wire_out_cluster_sb_BR_2_3, wire_out_cluster_sb_BR_1_3, wire_out_cluster_sb_BR_0_3 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_3, wire_out_cluster_sb_TL_2_3, wire_out_cluster_sb_TL_1_3, wire_out_cluster_sb_TL_0_3 } )
      , .outpads_0( outpads_right[0] )
      , .outpads_1( outpads_top[0] )
      , .sb_bottom_input( { wire_sb_bottom_input_11_4, wire_sb_bottom_input_10_4, wire_sb_bottom_input_9_4, wire_sb_bottom_input_8_4, wire_sb_bottom_input_7_4, wire_sb_bottom_input_6_4, wire_sb_bottom_input_5_4, wire_sb_bottom_input_4_4, wire_sb_bottom_input_3_4, wire_sb_bottom_input_2_4, wire_sb_bottom_input_1_4, wire_sb_bottom_input_0_4 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_4, wire_sb_bottom_output_10_4, wire_sb_bottom_output_9_4, wire_sb_bottom_output_8_4, wire_sb_bottom_output_7_4, wire_sb_bottom_output_6_4, wire_sb_bottom_output_5_4, wire_sb_bottom_output_4_4, wire_sb_bottom_output_3_4, wire_sb_bottom_output_2_4, wire_sb_bottom_output_1_4, wire_sb_bottom_output_0_4 } )
      , .sb_left_input( { wire_sb_left_input_11_3, wire_sb_left_input_10_3, wire_sb_left_input_9_3, wire_sb_left_input_8_3, wire_sb_left_input_7_3, wire_sb_left_input_6_3, wire_sb_left_input_5_3, wire_sb_left_input_4_3, wire_sb_left_input_3_3, wire_sb_left_input_2_3, wire_sb_left_input_1_3, wire_sb_left_input_0_3 } )
      , .sb_left_output( { wire_sb_left_output_11_3, wire_sb_left_output_10_3, wire_sb_left_output_9_3, wire_sb_left_output_8_3, wire_sb_left_output_7_3, wire_sb_left_output_6_3, wire_sb_left_output_5_3, wire_sb_left_output_4_3, wire_sb_left_output_3_3, wire_sb_left_output_2_3, wire_sb_left_output_1_3, wire_sb_left_output_0_3 } )
     );

TileInternal tile_I11(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[11] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_9, wire_in_cluster_sb_TL_14_9, wire_in_cluster_sb_TL_13_9, wire_in_cluster_sb_TL_12_9, wire_in_cluster_sb_TL_11_9, wire_in_cluster_sb_TL_10_9, wire_in_cluster_sb_TL_9_9, wire_in_cluster_sb_TL_8_9, wire_in_cluster_sb_TL_7_9, wire_in_cluster_sb_TL_6_9, wire_in_cluster_sb_TL_5_9, wire_in_cluster_sb_TL_4_9, wire_in_cluster_sb_TL_3_9, wire_in_cluster_sb_TL_2_9, wire_in_cluster_sb_TL_1_9, wire_in_cluster_sb_TL_0_9 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_4, wire_in_cluster_sb_BR_14_4, wire_in_cluster_sb_BR_13_4, wire_in_cluster_sb_BR_12_4, wire_in_cluster_sb_BR_11_4, wire_in_cluster_sb_BR_10_4, wire_in_cluster_sb_BR_9_4, wire_in_cluster_sb_BR_8_4, wire_in_cluster_sb_BR_7_4, wire_in_cluster_sb_BR_6_4, wire_in_cluster_sb_BR_5_4, wire_in_cluster_sb_BR_4_4, wire_in_cluster_sb_BR_3_4, wire_in_cluster_sb_BR_2_4, wire_in_cluster_sb_BR_1_4, wire_in_cluster_sb_BR_0_4 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_5, wire_in_cluster_sb_BL_14_5, wire_in_cluster_sb_BL_13_5, wire_in_cluster_sb_BL_12_5, wire_in_cluster_sb_BL_11_5, wire_in_cluster_sb_BL_10_5, wire_in_cluster_sb_BL_9_5, wire_in_cluster_sb_BL_8_5, wire_in_cluster_sb_BL_7_5, wire_in_cluster_sb_BL_6_5, wire_in_cluster_sb_BL_5_5, wire_in_cluster_sb_BL_4_5, wire_in_cluster_sb_BL_3_5, wire_in_cluster_sb_BL_2_5, wire_in_cluster_sb_BL_1_5, wire_in_cluster_sb_BL_0_5 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_8, wire_in_cluster_sb_BL_14_8, wire_in_cluster_sb_BL_13_8, wire_in_cluster_sb_BL_12_8, wire_in_cluster_sb_BL_11_8, wire_in_cluster_sb_BL_10_8, wire_in_cluster_sb_BL_9_8, wire_in_cluster_sb_BL_8_8, wire_in_cluster_sb_BL_7_8, wire_in_cluster_sb_BL_6_8, wire_in_cluster_sb_BL_5_8, wire_in_cluster_sb_BL_4_8, wire_in_cluster_sb_BL_3_8, wire_in_cluster_sb_BL_2_8, wire_in_cluster_sb_BL_1_8, wire_in_cluster_sb_BL_0_8 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_8, wire_in_cluster_sb_BR_14_8, wire_in_cluster_sb_BR_13_8, wire_in_cluster_sb_BR_12_8, wire_in_cluster_sb_BR_11_8, wire_in_cluster_sb_BR_10_8, wire_in_cluster_sb_BR_9_8, wire_in_cluster_sb_BR_8_8, wire_in_cluster_sb_BR_7_8, wire_in_cluster_sb_BR_6_8, wire_in_cluster_sb_BR_5_8, wire_in_cluster_sb_BR_4_8, wire_in_cluster_sb_BR_3_8, wire_in_cluster_sb_BR_2_8, wire_in_cluster_sb_BR_1_8, wire_in_cluster_sb_BR_0_8 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_8, wire_in_cluster_sb_TL_14_8, wire_in_cluster_sb_TL_13_8, wire_in_cluster_sb_TL_12_8, wire_in_cluster_sb_TL_11_8, wire_in_cluster_sb_TL_10_8, wire_in_cluster_sb_TL_9_8, wire_in_cluster_sb_TL_8_8, wire_in_cluster_sb_TL_7_8, wire_in_cluster_sb_TL_6_8, wire_in_cluster_sb_TL_5_8, wire_in_cluster_sb_TL_4_8, wire_in_cluster_sb_TL_3_8, wire_in_cluster_sb_TL_2_8, wire_in_cluster_sb_TL_1_8, wire_in_cluster_sb_TL_0_8 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_9, wire_out_cluster_sb_TL_2_9, wire_out_cluster_sb_TL_1_9, wire_out_cluster_sb_TL_0_9 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_4, wire_out_cluster_sb_BR_2_4, wire_out_cluster_sb_BR_1_4, wire_out_cluster_sb_BR_0_4 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_5, wire_out_cluster_sb_BL_2_5, wire_out_cluster_sb_BL_1_5, wire_out_cluster_sb_BL_0_5 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_8, wire_out_cluster_sb_BL_2_8, wire_out_cluster_sb_BL_1_8, wire_out_cluster_sb_BL_0_8 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_8, wire_out_cluster_sb_BR_2_8, wire_out_cluster_sb_BR_1_8, wire_out_cluster_sb_BR_0_8 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_8, wire_out_cluster_sb_TL_2_8, wire_out_cluster_sb_TL_1_8, wire_out_cluster_sb_TL_0_8 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_11, wire_sb_bottom_input_10_11, wire_sb_bottom_input_9_11, wire_sb_bottom_input_8_11, wire_sb_bottom_input_7_11, wire_sb_bottom_input_6_11, wire_sb_bottom_input_5_11, wire_sb_bottom_input_4_11, wire_sb_bottom_input_3_11, wire_sb_bottom_input_2_11, wire_sb_bottom_input_1_11, wire_sb_bottom_input_0_11 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_11, wire_sb_bottom_output_10_11, wire_sb_bottom_output_9_11, wire_sb_bottom_output_8_11, wire_sb_bottom_output_7_11, wire_sb_bottom_output_6_11, wire_sb_bottom_output_5_11, wire_sb_bottom_output_4_11, wire_sb_bottom_output_3_11, wire_sb_bottom_output_2_11, wire_sb_bottom_output_1_11, wire_sb_bottom_output_0_11 } )
      , .sb_left_input( { wire_sb_left_input_11_8, wire_sb_left_input_10_8, wire_sb_left_input_9_8, wire_sb_left_input_8_8, wire_sb_left_input_7_8, wire_sb_left_input_6_8, wire_sb_left_input_5_8, wire_sb_left_input_4_8, wire_sb_left_input_3_8, wire_sb_left_input_2_8, wire_sb_left_input_1_8, wire_sb_left_input_0_8 } )
      , .sb_left_output( { wire_sb_left_output_11_8, wire_sb_left_output_10_8, wire_sb_left_output_9_8, wire_sb_left_output_8_8, wire_sb_left_output_7_8, wire_sb_left_output_6_8, wire_sb_left_output_5_8, wire_sb_left_output_4_8, wire_sb_left_output_3_8, wire_sb_left_output_2_8, wire_sb_left_output_1_8, wire_sb_left_output_0_8 } )
      , .sb_right_input( { wire_sb_left_output_11_9, wire_sb_left_output_10_9, wire_sb_left_output_9_9, wire_sb_left_output_8_9, wire_sb_left_output_7_9, wire_sb_left_output_6_9, wire_sb_left_output_5_9, wire_sb_left_output_4_9, wire_sb_left_output_3_9, wire_sb_left_output_2_9, wire_sb_left_output_1_9, wire_sb_left_output_0_9 } )
      , .sb_right_output( { wire_sb_left_input_11_9, wire_sb_left_input_10_9, wire_sb_left_input_9_9, wire_sb_left_input_8_9, wire_sb_left_input_7_9, wire_sb_left_input_6_9, wire_sb_left_input_5_9, wire_sb_left_input_4_9, wire_sb_left_input_3_9, wire_sb_left_input_2_9, wire_sb_left_input_1_9, wire_sb_left_input_0_9 } )
      , .sb_top_input( { wire_sb_bottom_output_11_6, wire_sb_bottom_output_10_6, wire_sb_bottom_output_9_6, wire_sb_bottom_output_8_6, wire_sb_bottom_output_7_6, wire_sb_bottom_output_6_6, wire_sb_bottom_output_5_6, wire_sb_bottom_output_4_6, wire_sb_bottom_output_3_6, wire_sb_bottom_output_2_6, wire_sb_bottom_output_1_6, wire_sb_bottom_output_0_6 } )
      , .sb_top_output( { wire_sb_bottom_input_11_6, wire_sb_bottom_input_10_6, wire_sb_bottom_input_9_6, wire_sb_bottom_input_8_6, wire_sb_bottom_input_7_6, wire_sb_bottom_input_6_6, wire_sb_bottom_input_5_6, wire_sb_bottom_input_4_6, wire_sb_bottom_input_3_6, wire_sb_bottom_input_2_6, wire_sb_bottom_input_1_6, wire_sb_bottom_input_0_6 } )
     );

TileInternal tile_I12(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[12] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_10, wire_in_cluster_sb_TL_14_10, wire_in_cluster_sb_TL_13_10, wire_in_cluster_sb_TL_12_10, wire_in_cluster_sb_TL_11_10, wire_in_cluster_sb_TL_10_10, wire_in_cluster_sb_TL_9_10, wire_in_cluster_sb_TL_8_10, wire_in_cluster_sb_TL_7_10, wire_in_cluster_sb_TL_6_10, wire_in_cluster_sb_TL_5_10, wire_in_cluster_sb_TL_4_10, wire_in_cluster_sb_TL_3_10, wire_in_cluster_sb_TL_2_10, wire_in_cluster_sb_TL_1_10, wire_in_cluster_sb_TL_0_10 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_5, wire_in_cluster_sb_BR_14_5, wire_in_cluster_sb_BR_13_5, wire_in_cluster_sb_BR_12_5, wire_in_cluster_sb_BR_11_5, wire_in_cluster_sb_BR_10_5, wire_in_cluster_sb_BR_9_5, wire_in_cluster_sb_BR_8_5, wire_in_cluster_sb_BR_7_5, wire_in_cluster_sb_BR_6_5, wire_in_cluster_sb_BR_5_5, wire_in_cluster_sb_BR_4_5, wire_in_cluster_sb_BR_3_5, wire_in_cluster_sb_BR_2_5, wire_in_cluster_sb_BR_1_5, wire_in_cluster_sb_BR_0_5 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_6, wire_in_cluster_sb_BL_14_6, wire_in_cluster_sb_BL_13_6, wire_in_cluster_sb_BL_12_6, wire_in_cluster_sb_BL_11_6, wire_in_cluster_sb_BL_10_6, wire_in_cluster_sb_BL_9_6, wire_in_cluster_sb_BL_8_6, wire_in_cluster_sb_BL_7_6, wire_in_cluster_sb_BL_6_6, wire_in_cluster_sb_BL_5_6, wire_in_cluster_sb_BL_4_6, wire_in_cluster_sb_BL_3_6, wire_in_cluster_sb_BL_2_6, wire_in_cluster_sb_BL_1_6, wire_in_cluster_sb_BL_0_6 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_9, wire_in_cluster_sb_BL_14_9, wire_in_cluster_sb_BL_13_9, wire_in_cluster_sb_BL_12_9, wire_in_cluster_sb_BL_11_9, wire_in_cluster_sb_BL_10_9, wire_in_cluster_sb_BL_9_9, wire_in_cluster_sb_BL_8_9, wire_in_cluster_sb_BL_7_9, wire_in_cluster_sb_BL_6_9, wire_in_cluster_sb_BL_5_9, wire_in_cluster_sb_BL_4_9, wire_in_cluster_sb_BL_3_9, wire_in_cluster_sb_BL_2_9, wire_in_cluster_sb_BL_1_9, wire_in_cluster_sb_BL_0_9 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_9, wire_in_cluster_sb_BR_14_9, wire_in_cluster_sb_BR_13_9, wire_in_cluster_sb_BR_12_9, wire_in_cluster_sb_BR_11_9, wire_in_cluster_sb_BR_10_9, wire_in_cluster_sb_BR_9_9, wire_in_cluster_sb_BR_8_9, wire_in_cluster_sb_BR_7_9, wire_in_cluster_sb_BR_6_9, wire_in_cluster_sb_BR_5_9, wire_in_cluster_sb_BR_4_9, wire_in_cluster_sb_BR_3_9, wire_in_cluster_sb_BR_2_9, wire_in_cluster_sb_BR_1_9, wire_in_cluster_sb_BR_0_9 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_9, wire_in_cluster_sb_TL_14_9, wire_in_cluster_sb_TL_13_9, wire_in_cluster_sb_TL_12_9, wire_in_cluster_sb_TL_11_9, wire_in_cluster_sb_TL_10_9, wire_in_cluster_sb_TL_9_9, wire_in_cluster_sb_TL_8_9, wire_in_cluster_sb_TL_7_9, wire_in_cluster_sb_TL_6_9, wire_in_cluster_sb_TL_5_9, wire_in_cluster_sb_TL_4_9, wire_in_cluster_sb_TL_3_9, wire_in_cluster_sb_TL_2_9, wire_in_cluster_sb_TL_1_9, wire_in_cluster_sb_TL_0_9 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_10, wire_out_cluster_sb_TL_2_10, wire_out_cluster_sb_TL_1_10, wire_out_cluster_sb_TL_0_10 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_5, wire_out_cluster_sb_BR_2_5, wire_out_cluster_sb_BR_1_5, wire_out_cluster_sb_BR_0_5 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_6, wire_out_cluster_sb_BL_2_6, wire_out_cluster_sb_BL_1_6, wire_out_cluster_sb_BL_0_6 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_9, wire_out_cluster_sb_BL_2_9, wire_out_cluster_sb_BL_1_9, wire_out_cluster_sb_BL_0_9 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_9, wire_out_cluster_sb_BR_2_9, wire_out_cluster_sb_BR_1_9, wire_out_cluster_sb_BR_0_9 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_9, wire_out_cluster_sb_TL_2_9, wire_out_cluster_sb_TL_1_9, wire_out_cluster_sb_TL_0_9 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_12, wire_sb_bottom_input_10_12, wire_sb_bottom_input_9_12, wire_sb_bottom_input_8_12, wire_sb_bottom_input_7_12, wire_sb_bottom_input_6_12, wire_sb_bottom_input_5_12, wire_sb_bottom_input_4_12, wire_sb_bottom_input_3_12, wire_sb_bottom_input_2_12, wire_sb_bottom_input_1_12, wire_sb_bottom_input_0_12 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_12, wire_sb_bottom_output_10_12, wire_sb_bottom_output_9_12, wire_sb_bottom_output_8_12, wire_sb_bottom_output_7_12, wire_sb_bottom_output_6_12, wire_sb_bottom_output_5_12, wire_sb_bottom_output_4_12, wire_sb_bottom_output_3_12, wire_sb_bottom_output_2_12, wire_sb_bottom_output_1_12, wire_sb_bottom_output_0_12 } )
      , .sb_left_input( { wire_sb_left_input_11_9, wire_sb_left_input_10_9, wire_sb_left_input_9_9, wire_sb_left_input_8_9, wire_sb_left_input_7_9, wire_sb_left_input_6_9, wire_sb_left_input_5_9, wire_sb_left_input_4_9, wire_sb_left_input_3_9, wire_sb_left_input_2_9, wire_sb_left_input_1_9, wire_sb_left_input_0_9 } )
      , .sb_left_output( { wire_sb_left_output_11_9, wire_sb_left_output_10_9, wire_sb_left_output_9_9, wire_sb_left_output_8_9, wire_sb_left_output_7_9, wire_sb_left_output_6_9, wire_sb_left_output_5_9, wire_sb_left_output_4_9, wire_sb_left_output_3_9, wire_sb_left_output_2_9, wire_sb_left_output_1_9, wire_sb_left_output_0_9 } )
      , .sb_right_input( { wire_sb_left_output_11_10, wire_sb_left_output_10_10, wire_sb_left_output_9_10, wire_sb_left_output_8_10, wire_sb_left_output_7_10, wire_sb_left_output_6_10, wire_sb_left_output_5_10, wire_sb_left_output_4_10, wire_sb_left_output_3_10, wire_sb_left_output_2_10, wire_sb_left_output_1_10, wire_sb_left_output_0_10 } )
      , .sb_right_output( { wire_sb_left_input_11_10, wire_sb_left_input_10_10, wire_sb_left_input_9_10, wire_sb_left_input_8_10, wire_sb_left_input_7_10, wire_sb_left_input_6_10, wire_sb_left_input_5_10, wire_sb_left_input_4_10, wire_sb_left_input_3_10, wire_sb_left_input_2_10, wire_sb_left_input_1_10, wire_sb_left_input_0_10 } )
      , .sb_top_input( { wire_sb_bottom_output_11_7, wire_sb_bottom_output_10_7, wire_sb_bottom_output_9_7, wire_sb_bottom_output_8_7, wire_sb_bottom_output_7_7, wire_sb_bottom_output_6_7, wire_sb_bottom_output_5_7, wire_sb_bottom_output_4_7, wire_sb_bottom_output_3_7, wire_sb_bottom_output_2_7, wire_sb_bottom_output_1_7, wire_sb_bottom_output_0_7 } )
      , .sb_top_output( { wire_sb_bottom_input_11_7, wire_sb_bottom_input_10_7, wire_sb_bottom_input_9_7, wire_sb_bottom_input_8_7, wire_sb_bottom_input_7_7, wire_sb_bottom_input_6_7, wire_sb_bottom_input_5_7, wire_sb_bottom_input_4_7, wire_sb_bottom_input_3_7, wire_sb_bottom_input_2_7, wire_sb_bottom_input_1_7, wire_sb_bottom_input_0_7 } )
     );

TileInternal tile_I13(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[13] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_11, wire_in_cluster_sb_TL_14_11, wire_in_cluster_sb_TL_13_11, wire_in_cluster_sb_TL_12_11, wire_in_cluster_sb_TL_11_11, wire_in_cluster_sb_TL_10_11, wire_in_cluster_sb_TL_9_11, wire_in_cluster_sb_TL_8_11, wire_in_cluster_sb_TL_7_11, wire_in_cluster_sb_TL_6_11, wire_in_cluster_sb_TL_5_11, wire_in_cluster_sb_TL_4_11, wire_in_cluster_sb_TL_3_11, wire_in_cluster_sb_TL_2_11, wire_in_cluster_sb_TL_1_11, wire_in_cluster_sb_TL_0_11 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_6, wire_in_cluster_sb_BR_14_6, wire_in_cluster_sb_BR_13_6, wire_in_cluster_sb_BR_12_6, wire_in_cluster_sb_BR_11_6, wire_in_cluster_sb_BR_10_6, wire_in_cluster_sb_BR_9_6, wire_in_cluster_sb_BR_8_6, wire_in_cluster_sb_BR_7_6, wire_in_cluster_sb_BR_6_6, wire_in_cluster_sb_BR_5_6, wire_in_cluster_sb_BR_4_6, wire_in_cluster_sb_BR_3_6, wire_in_cluster_sb_BR_2_6, wire_in_cluster_sb_BR_1_6, wire_in_cluster_sb_BR_0_6 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_7, wire_in_cluster_sb_BL_14_7, wire_in_cluster_sb_BL_13_7, wire_in_cluster_sb_BL_12_7, wire_in_cluster_sb_BL_11_7, wire_in_cluster_sb_BL_10_7, wire_in_cluster_sb_BL_9_7, wire_in_cluster_sb_BL_8_7, wire_in_cluster_sb_BL_7_7, wire_in_cluster_sb_BL_6_7, wire_in_cluster_sb_BL_5_7, wire_in_cluster_sb_BL_4_7, wire_in_cluster_sb_BL_3_7, wire_in_cluster_sb_BL_2_7, wire_in_cluster_sb_BL_1_7, wire_in_cluster_sb_BL_0_7 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_10, wire_in_cluster_sb_BL_14_10, wire_in_cluster_sb_BL_13_10, wire_in_cluster_sb_BL_12_10, wire_in_cluster_sb_BL_11_10, wire_in_cluster_sb_BL_10_10, wire_in_cluster_sb_BL_9_10, wire_in_cluster_sb_BL_8_10, wire_in_cluster_sb_BL_7_10, wire_in_cluster_sb_BL_6_10, wire_in_cluster_sb_BL_5_10, wire_in_cluster_sb_BL_4_10, wire_in_cluster_sb_BL_3_10, wire_in_cluster_sb_BL_2_10, wire_in_cluster_sb_BL_1_10, wire_in_cluster_sb_BL_0_10 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_10, wire_in_cluster_sb_BR_14_10, wire_in_cluster_sb_BR_13_10, wire_in_cluster_sb_BR_12_10, wire_in_cluster_sb_BR_11_10, wire_in_cluster_sb_BR_10_10, wire_in_cluster_sb_BR_9_10, wire_in_cluster_sb_BR_8_10, wire_in_cluster_sb_BR_7_10, wire_in_cluster_sb_BR_6_10, wire_in_cluster_sb_BR_5_10, wire_in_cluster_sb_BR_4_10, wire_in_cluster_sb_BR_3_10, wire_in_cluster_sb_BR_2_10, wire_in_cluster_sb_BR_1_10, wire_in_cluster_sb_BR_0_10 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_10, wire_in_cluster_sb_TL_14_10, wire_in_cluster_sb_TL_13_10, wire_in_cluster_sb_TL_12_10, wire_in_cluster_sb_TL_11_10, wire_in_cluster_sb_TL_10_10, wire_in_cluster_sb_TL_9_10, wire_in_cluster_sb_TL_8_10, wire_in_cluster_sb_TL_7_10, wire_in_cluster_sb_TL_6_10, wire_in_cluster_sb_TL_5_10, wire_in_cluster_sb_TL_4_10, wire_in_cluster_sb_TL_3_10, wire_in_cluster_sb_TL_2_10, wire_in_cluster_sb_TL_1_10, wire_in_cluster_sb_TL_0_10 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_11, wire_out_cluster_sb_TL_2_11, wire_out_cluster_sb_TL_1_11, wire_out_cluster_sb_TL_0_11 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_6, wire_out_cluster_sb_BR_2_6, wire_out_cluster_sb_BR_1_6, wire_out_cluster_sb_BR_0_6 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_7, wire_out_cluster_sb_BL_2_7, wire_out_cluster_sb_BL_1_7, wire_out_cluster_sb_BL_0_7 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_10, wire_out_cluster_sb_BL_2_10, wire_out_cluster_sb_BL_1_10, wire_out_cluster_sb_BL_0_10 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_10, wire_out_cluster_sb_BR_2_10, wire_out_cluster_sb_BR_1_10, wire_out_cluster_sb_BR_0_10 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_10, wire_out_cluster_sb_TL_2_10, wire_out_cluster_sb_TL_1_10, wire_out_cluster_sb_TL_0_10 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_13, wire_sb_bottom_input_10_13, wire_sb_bottom_input_9_13, wire_sb_bottom_input_8_13, wire_sb_bottom_input_7_13, wire_sb_bottom_input_6_13, wire_sb_bottom_input_5_13, wire_sb_bottom_input_4_13, wire_sb_bottom_input_3_13, wire_sb_bottom_input_2_13, wire_sb_bottom_input_1_13, wire_sb_bottom_input_0_13 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_13, wire_sb_bottom_output_10_13, wire_sb_bottom_output_9_13, wire_sb_bottom_output_8_13, wire_sb_bottom_output_7_13, wire_sb_bottom_output_6_13, wire_sb_bottom_output_5_13, wire_sb_bottom_output_4_13, wire_sb_bottom_output_3_13, wire_sb_bottom_output_2_13, wire_sb_bottom_output_1_13, wire_sb_bottom_output_0_13 } )
      , .sb_left_input( { wire_sb_left_input_11_10, wire_sb_left_input_10_10, wire_sb_left_input_9_10, wire_sb_left_input_8_10, wire_sb_left_input_7_10, wire_sb_left_input_6_10, wire_sb_left_input_5_10, wire_sb_left_input_4_10, wire_sb_left_input_3_10, wire_sb_left_input_2_10, wire_sb_left_input_1_10, wire_sb_left_input_0_10 } )
      , .sb_left_output( { wire_sb_left_output_11_10, wire_sb_left_output_10_10, wire_sb_left_output_9_10, wire_sb_left_output_8_10, wire_sb_left_output_7_10, wire_sb_left_output_6_10, wire_sb_left_output_5_10, wire_sb_left_output_4_10, wire_sb_left_output_3_10, wire_sb_left_output_2_10, wire_sb_left_output_1_10, wire_sb_left_output_0_10 } )
      , .sb_right_input( { wire_sb_left_output_11_11, wire_sb_left_output_10_11, wire_sb_left_output_9_11, wire_sb_left_output_8_11, wire_sb_left_output_7_11, wire_sb_left_output_6_11, wire_sb_left_output_5_11, wire_sb_left_output_4_11, wire_sb_left_output_3_11, wire_sb_left_output_2_11, wire_sb_left_output_1_11, wire_sb_left_output_0_11 } )
      , .sb_right_output( { wire_sb_left_input_11_11, wire_sb_left_input_10_11, wire_sb_left_input_9_11, wire_sb_left_input_8_11, wire_sb_left_input_7_11, wire_sb_left_input_6_11, wire_sb_left_input_5_11, wire_sb_left_input_4_11, wire_sb_left_input_3_11, wire_sb_left_input_2_11, wire_sb_left_input_1_11, wire_sb_left_input_0_11 } )
      , .sb_top_input( { wire_sb_bottom_output_11_8, wire_sb_bottom_output_10_8, wire_sb_bottom_output_9_8, wire_sb_bottom_output_8_8, wire_sb_bottom_output_7_8, wire_sb_bottom_output_6_8, wire_sb_bottom_output_5_8, wire_sb_bottom_output_4_8, wire_sb_bottom_output_3_8, wire_sb_bottom_output_2_8, wire_sb_bottom_output_1_8, wire_sb_bottom_output_0_8 } )
      , .sb_top_output( { wire_sb_bottom_input_11_8, wire_sb_bottom_input_10_8, wire_sb_bottom_input_9_8, wire_sb_bottom_input_8_8, wire_sb_bottom_input_7_8, wire_sb_bottom_input_6_8, wire_sb_bottom_input_5_8, wire_sb_bottom_input_4_8, wire_sb_bottom_input_3_8, wire_sb_bottom_input_2_8, wire_sb_bottom_input_1_8, wire_sb_bottom_input_0_8 } )
     );

TileInternal tile_I16(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[16] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_13, wire_in_cluster_sb_TL_14_13, wire_in_cluster_sb_TL_13_13, wire_in_cluster_sb_TL_12_13, wire_in_cluster_sb_TL_11_13, wire_in_cluster_sb_TL_10_13, wire_in_cluster_sb_TL_9_13, wire_in_cluster_sb_TL_8_13, wire_in_cluster_sb_TL_7_13, wire_in_cluster_sb_TL_6_13, wire_in_cluster_sb_TL_5_13, wire_in_cluster_sb_TL_4_13, wire_in_cluster_sb_TL_3_13, wire_in_cluster_sb_TL_2_13, wire_in_cluster_sb_TL_1_13, wire_in_cluster_sb_TL_0_13 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_8, wire_in_cluster_sb_BR_14_8, wire_in_cluster_sb_BR_13_8, wire_in_cluster_sb_BR_12_8, wire_in_cluster_sb_BR_11_8, wire_in_cluster_sb_BR_10_8, wire_in_cluster_sb_BR_9_8, wire_in_cluster_sb_BR_8_8, wire_in_cluster_sb_BR_7_8, wire_in_cluster_sb_BR_6_8, wire_in_cluster_sb_BR_5_8, wire_in_cluster_sb_BR_4_8, wire_in_cluster_sb_BR_3_8, wire_in_cluster_sb_BR_2_8, wire_in_cluster_sb_BR_1_8, wire_in_cluster_sb_BR_0_8 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_9, wire_in_cluster_sb_BL_14_9, wire_in_cluster_sb_BL_13_9, wire_in_cluster_sb_BL_12_9, wire_in_cluster_sb_BL_11_9, wire_in_cluster_sb_BL_10_9, wire_in_cluster_sb_BL_9_9, wire_in_cluster_sb_BL_8_9, wire_in_cluster_sb_BL_7_9, wire_in_cluster_sb_BL_6_9, wire_in_cluster_sb_BL_5_9, wire_in_cluster_sb_BL_4_9, wire_in_cluster_sb_BL_3_9, wire_in_cluster_sb_BL_2_9, wire_in_cluster_sb_BL_1_9, wire_in_cluster_sb_BL_0_9 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_12, wire_in_cluster_sb_BL_14_12, wire_in_cluster_sb_BL_13_12, wire_in_cluster_sb_BL_12_12, wire_in_cluster_sb_BL_11_12, wire_in_cluster_sb_BL_10_12, wire_in_cluster_sb_BL_9_12, wire_in_cluster_sb_BL_8_12, wire_in_cluster_sb_BL_7_12, wire_in_cluster_sb_BL_6_12, wire_in_cluster_sb_BL_5_12, wire_in_cluster_sb_BL_4_12, wire_in_cluster_sb_BL_3_12, wire_in_cluster_sb_BL_2_12, wire_in_cluster_sb_BL_1_12, wire_in_cluster_sb_BL_0_12 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_12, wire_in_cluster_sb_BR_14_12, wire_in_cluster_sb_BR_13_12, wire_in_cluster_sb_BR_12_12, wire_in_cluster_sb_BR_11_12, wire_in_cluster_sb_BR_10_12, wire_in_cluster_sb_BR_9_12, wire_in_cluster_sb_BR_8_12, wire_in_cluster_sb_BR_7_12, wire_in_cluster_sb_BR_6_12, wire_in_cluster_sb_BR_5_12, wire_in_cluster_sb_BR_4_12, wire_in_cluster_sb_BR_3_12, wire_in_cluster_sb_BR_2_12, wire_in_cluster_sb_BR_1_12, wire_in_cluster_sb_BR_0_12 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_12, wire_in_cluster_sb_TL_14_12, wire_in_cluster_sb_TL_13_12, wire_in_cluster_sb_TL_12_12, wire_in_cluster_sb_TL_11_12, wire_in_cluster_sb_TL_10_12, wire_in_cluster_sb_TL_9_12, wire_in_cluster_sb_TL_8_12, wire_in_cluster_sb_TL_7_12, wire_in_cluster_sb_TL_6_12, wire_in_cluster_sb_TL_5_12, wire_in_cluster_sb_TL_4_12, wire_in_cluster_sb_TL_3_12, wire_in_cluster_sb_TL_2_12, wire_in_cluster_sb_TL_1_12, wire_in_cluster_sb_TL_0_12 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_13, wire_out_cluster_sb_TL_2_13, wire_out_cluster_sb_TL_1_13, wire_out_cluster_sb_TL_0_13 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_8, wire_out_cluster_sb_BR_2_8, wire_out_cluster_sb_BR_1_8, wire_out_cluster_sb_BR_0_8 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_9, wire_out_cluster_sb_BL_2_9, wire_out_cluster_sb_BL_1_9, wire_out_cluster_sb_BL_0_9 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_12, wire_out_cluster_sb_BL_2_12, wire_out_cluster_sb_BL_1_12, wire_out_cluster_sb_BL_0_12 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_12, wire_out_cluster_sb_BR_2_12, wire_out_cluster_sb_BR_1_12, wire_out_cluster_sb_BR_0_12 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_12, wire_out_cluster_sb_TL_2_12, wire_out_cluster_sb_TL_1_12, wire_out_cluster_sb_TL_0_12 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_16, wire_sb_bottom_input_10_16, wire_sb_bottom_input_9_16, wire_sb_bottom_input_8_16, wire_sb_bottom_input_7_16, wire_sb_bottom_input_6_16, wire_sb_bottom_input_5_16, wire_sb_bottom_input_4_16, wire_sb_bottom_input_3_16, wire_sb_bottom_input_2_16, wire_sb_bottom_input_1_16, wire_sb_bottom_input_0_16 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_16, wire_sb_bottom_output_10_16, wire_sb_bottom_output_9_16, wire_sb_bottom_output_8_16, wire_sb_bottom_output_7_16, wire_sb_bottom_output_6_16, wire_sb_bottom_output_5_16, wire_sb_bottom_output_4_16, wire_sb_bottom_output_3_16, wire_sb_bottom_output_2_16, wire_sb_bottom_output_1_16, wire_sb_bottom_output_0_16 } )
      , .sb_left_input( { wire_sb_left_input_11_12, wire_sb_left_input_10_12, wire_sb_left_input_9_12, wire_sb_left_input_8_12, wire_sb_left_input_7_12, wire_sb_left_input_6_12, wire_sb_left_input_5_12, wire_sb_left_input_4_12, wire_sb_left_input_3_12, wire_sb_left_input_2_12, wire_sb_left_input_1_12, wire_sb_left_input_0_12 } )
      , .sb_left_output( { wire_sb_left_output_11_12, wire_sb_left_output_10_12, wire_sb_left_output_9_12, wire_sb_left_output_8_12, wire_sb_left_output_7_12, wire_sb_left_output_6_12, wire_sb_left_output_5_12, wire_sb_left_output_4_12, wire_sb_left_output_3_12, wire_sb_left_output_2_12, wire_sb_left_output_1_12, wire_sb_left_output_0_12 } )
      , .sb_right_input( { wire_sb_left_output_11_13, wire_sb_left_output_10_13, wire_sb_left_output_9_13, wire_sb_left_output_8_13, wire_sb_left_output_7_13, wire_sb_left_output_6_13, wire_sb_left_output_5_13, wire_sb_left_output_4_13, wire_sb_left_output_3_13, wire_sb_left_output_2_13, wire_sb_left_output_1_13, wire_sb_left_output_0_13 } )
      , .sb_right_output( { wire_sb_left_input_11_13, wire_sb_left_input_10_13, wire_sb_left_input_9_13, wire_sb_left_input_8_13, wire_sb_left_input_7_13, wire_sb_left_input_6_13, wire_sb_left_input_5_13, wire_sb_left_input_4_13, wire_sb_left_input_3_13, wire_sb_left_input_2_13, wire_sb_left_input_1_13, wire_sb_left_input_0_13 } )
      , .sb_top_input( { wire_sb_bottom_output_11_11, wire_sb_bottom_output_10_11, wire_sb_bottom_output_9_11, wire_sb_bottom_output_8_11, wire_sb_bottom_output_7_11, wire_sb_bottom_output_6_11, wire_sb_bottom_output_5_11, wire_sb_bottom_output_4_11, wire_sb_bottom_output_3_11, wire_sb_bottom_output_2_11, wire_sb_bottom_output_1_11, wire_sb_bottom_output_0_11 } )
      , .sb_top_output( { wire_sb_bottom_input_11_11, wire_sb_bottom_input_10_11, wire_sb_bottom_input_9_11, wire_sb_bottom_input_8_11, wire_sb_bottom_input_7_11, wire_sb_bottom_input_6_11, wire_sb_bottom_input_5_11, wire_sb_bottom_input_4_11, wire_sb_bottom_input_3_11, wire_sb_bottom_input_2_11, wire_sb_bottom_input_1_11, wire_sb_bottom_input_0_11 } )
     );

TileInternal tile_I17(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[17] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_14, wire_in_cluster_sb_TL_14_14, wire_in_cluster_sb_TL_13_14, wire_in_cluster_sb_TL_12_14, wire_in_cluster_sb_TL_11_14, wire_in_cluster_sb_TL_10_14, wire_in_cluster_sb_TL_9_14, wire_in_cluster_sb_TL_8_14, wire_in_cluster_sb_TL_7_14, wire_in_cluster_sb_TL_6_14, wire_in_cluster_sb_TL_5_14, wire_in_cluster_sb_TL_4_14, wire_in_cluster_sb_TL_3_14, wire_in_cluster_sb_TL_2_14, wire_in_cluster_sb_TL_1_14, wire_in_cluster_sb_TL_0_14 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_9, wire_in_cluster_sb_BR_14_9, wire_in_cluster_sb_BR_13_9, wire_in_cluster_sb_BR_12_9, wire_in_cluster_sb_BR_11_9, wire_in_cluster_sb_BR_10_9, wire_in_cluster_sb_BR_9_9, wire_in_cluster_sb_BR_8_9, wire_in_cluster_sb_BR_7_9, wire_in_cluster_sb_BR_6_9, wire_in_cluster_sb_BR_5_9, wire_in_cluster_sb_BR_4_9, wire_in_cluster_sb_BR_3_9, wire_in_cluster_sb_BR_2_9, wire_in_cluster_sb_BR_1_9, wire_in_cluster_sb_BR_0_9 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_10, wire_in_cluster_sb_BL_14_10, wire_in_cluster_sb_BL_13_10, wire_in_cluster_sb_BL_12_10, wire_in_cluster_sb_BL_11_10, wire_in_cluster_sb_BL_10_10, wire_in_cluster_sb_BL_9_10, wire_in_cluster_sb_BL_8_10, wire_in_cluster_sb_BL_7_10, wire_in_cluster_sb_BL_6_10, wire_in_cluster_sb_BL_5_10, wire_in_cluster_sb_BL_4_10, wire_in_cluster_sb_BL_3_10, wire_in_cluster_sb_BL_2_10, wire_in_cluster_sb_BL_1_10, wire_in_cluster_sb_BL_0_10 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_13, wire_in_cluster_sb_BL_14_13, wire_in_cluster_sb_BL_13_13, wire_in_cluster_sb_BL_12_13, wire_in_cluster_sb_BL_11_13, wire_in_cluster_sb_BL_10_13, wire_in_cluster_sb_BL_9_13, wire_in_cluster_sb_BL_8_13, wire_in_cluster_sb_BL_7_13, wire_in_cluster_sb_BL_6_13, wire_in_cluster_sb_BL_5_13, wire_in_cluster_sb_BL_4_13, wire_in_cluster_sb_BL_3_13, wire_in_cluster_sb_BL_2_13, wire_in_cluster_sb_BL_1_13, wire_in_cluster_sb_BL_0_13 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_13, wire_in_cluster_sb_BR_14_13, wire_in_cluster_sb_BR_13_13, wire_in_cluster_sb_BR_12_13, wire_in_cluster_sb_BR_11_13, wire_in_cluster_sb_BR_10_13, wire_in_cluster_sb_BR_9_13, wire_in_cluster_sb_BR_8_13, wire_in_cluster_sb_BR_7_13, wire_in_cluster_sb_BR_6_13, wire_in_cluster_sb_BR_5_13, wire_in_cluster_sb_BR_4_13, wire_in_cluster_sb_BR_3_13, wire_in_cluster_sb_BR_2_13, wire_in_cluster_sb_BR_1_13, wire_in_cluster_sb_BR_0_13 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_13, wire_in_cluster_sb_TL_14_13, wire_in_cluster_sb_TL_13_13, wire_in_cluster_sb_TL_12_13, wire_in_cluster_sb_TL_11_13, wire_in_cluster_sb_TL_10_13, wire_in_cluster_sb_TL_9_13, wire_in_cluster_sb_TL_8_13, wire_in_cluster_sb_TL_7_13, wire_in_cluster_sb_TL_6_13, wire_in_cluster_sb_TL_5_13, wire_in_cluster_sb_TL_4_13, wire_in_cluster_sb_TL_3_13, wire_in_cluster_sb_TL_2_13, wire_in_cluster_sb_TL_1_13, wire_in_cluster_sb_TL_0_13 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_14, wire_out_cluster_sb_TL_2_14, wire_out_cluster_sb_TL_1_14, wire_out_cluster_sb_TL_0_14 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_9, wire_out_cluster_sb_BR_2_9, wire_out_cluster_sb_BR_1_9, wire_out_cluster_sb_BR_0_9 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_10, wire_out_cluster_sb_BL_2_10, wire_out_cluster_sb_BL_1_10, wire_out_cluster_sb_BL_0_10 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_13, wire_out_cluster_sb_BL_2_13, wire_out_cluster_sb_BL_1_13, wire_out_cluster_sb_BL_0_13 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_13, wire_out_cluster_sb_BR_2_13, wire_out_cluster_sb_BR_1_13, wire_out_cluster_sb_BR_0_13 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_13, wire_out_cluster_sb_TL_2_13, wire_out_cluster_sb_TL_1_13, wire_out_cluster_sb_TL_0_13 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_17, wire_sb_bottom_input_10_17, wire_sb_bottom_input_9_17, wire_sb_bottom_input_8_17, wire_sb_bottom_input_7_17, wire_sb_bottom_input_6_17, wire_sb_bottom_input_5_17, wire_sb_bottom_input_4_17, wire_sb_bottom_input_3_17, wire_sb_bottom_input_2_17, wire_sb_bottom_input_1_17, wire_sb_bottom_input_0_17 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_17, wire_sb_bottom_output_10_17, wire_sb_bottom_output_9_17, wire_sb_bottom_output_8_17, wire_sb_bottom_output_7_17, wire_sb_bottom_output_6_17, wire_sb_bottom_output_5_17, wire_sb_bottom_output_4_17, wire_sb_bottom_output_3_17, wire_sb_bottom_output_2_17, wire_sb_bottom_output_1_17, wire_sb_bottom_output_0_17 } )
      , .sb_left_input( { wire_sb_left_input_11_13, wire_sb_left_input_10_13, wire_sb_left_input_9_13, wire_sb_left_input_8_13, wire_sb_left_input_7_13, wire_sb_left_input_6_13, wire_sb_left_input_5_13, wire_sb_left_input_4_13, wire_sb_left_input_3_13, wire_sb_left_input_2_13, wire_sb_left_input_1_13, wire_sb_left_input_0_13 } )
      , .sb_left_output( { wire_sb_left_output_11_13, wire_sb_left_output_10_13, wire_sb_left_output_9_13, wire_sb_left_output_8_13, wire_sb_left_output_7_13, wire_sb_left_output_6_13, wire_sb_left_output_5_13, wire_sb_left_output_4_13, wire_sb_left_output_3_13, wire_sb_left_output_2_13, wire_sb_left_output_1_13, wire_sb_left_output_0_13 } )
      , .sb_right_input( { wire_sb_left_output_11_14, wire_sb_left_output_10_14, wire_sb_left_output_9_14, wire_sb_left_output_8_14, wire_sb_left_output_7_14, wire_sb_left_output_6_14, wire_sb_left_output_5_14, wire_sb_left_output_4_14, wire_sb_left_output_3_14, wire_sb_left_output_2_14, wire_sb_left_output_1_14, wire_sb_left_output_0_14 } )
      , .sb_right_output( { wire_sb_left_input_11_14, wire_sb_left_input_10_14, wire_sb_left_input_9_14, wire_sb_left_input_8_14, wire_sb_left_input_7_14, wire_sb_left_input_6_14, wire_sb_left_input_5_14, wire_sb_left_input_4_14, wire_sb_left_input_3_14, wire_sb_left_input_2_14, wire_sb_left_input_1_14, wire_sb_left_input_0_14 } )
      , .sb_top_input( { wire_sb_bottom_output_11_12, wire_sb_bottom_output_10_12, wire_sb_bottom_output_9_12, wire_sb_bottom_output_8_12, wire_sb_bottom_output_7_12, wire_sb_bottom_output_6_12, wire_sb_bottom_output_5_12, wire_sb_bottom_output_4_12, wire_sb_bottom_output_3_12, wire_sb_bottom_output_2_12, wire_sb_bottom_output_1_12, wire_sb_bottom_output_0_12 } )
      , .sb_top_output( { wire_sb_bottom_input_11_12, wire_sb_bottom_input_10_12, wire_sb_bottom_input_9_12, wire_sb_bottom_input_8_12, wire_sb_bottom_input_7_12, wire_sb_bottom_input_6_12, wire_sb_bottom_input_5_12, wire_sb_bottom_input_4_12, wire_sb_bottom_input_3_12, wire_sb_bottom_input_2_12, wire_sb_bottom_input_1_12, wire_sb_bottom_input_0_12 } )
     );

TileInternal tile_I18(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[18] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_15, wire_in_cluster_sb_TL_14_15, wire_in_cluster_sb_TL_13_15, wire_in_cluster_sb_TL_12_15, wire_in_cluster_sb_TL_11_15, wire_in_cluster_sb_TL_10_15, wire_in_cluster_sb_TL_9_15, wire_in_cluster_sb_TL_8_15, wire_in_cluster_sb_TL_7_15, wire_in_cluster_sb_TL_6_15, wire_in_cluster_sb_TL_5_15, wire_in_cluster_sb_TL_4_15, wire_in_cluster_sb_TL_3_15, wire_in_cluster_sb_TL_2_15, wire_in_cluster_sb_TL_1_15, wire_in_cluster_sb_TL_0_15 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_10, wire_in_cluster_sb_BR_14_10, wire_in_cluster_sb_BR_13_10, wire_in_cluster_sb_BR_12_10, wire_in_cluster_sb_BR_11_10, wire_in_cluster_sb_BR_10_10, wire_in_cluster_sb_BR_9_10, wire_in_cluster_sb_BR_8_10, wire_in_cluster_sb_BR_7_10, wire_in_cluster_sb_BR_6_10, wire_in_cluster_sb_BR_5_10, wire_in_cluster_sb_BR_4_10, wire_in_cluster_sb_BR_3_10, wire_in_cluster_sb_BR_2_10, wire_in_cluster_sb_BR_1_10, wire_in_cluster_sb_BR_0_10 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_11, wire_in_cluster_sb_BL_14_11, wire_in_cluster_sb_BL_13_11, wire_in_cluster_sb_BL_12_11, wire_in_cluster_sb_BL_11_11, wire_in_cluster_sb_BL_10_11, wire_in_cluster_sb_BL_9_11, wire_in_cluster_sb_BL_8_11, wire_in_cluster_sb_BL_7_11, wire_in_cluster_sb_BL_6_11, wire_in_cluster_sb_BL_5_11, wire_in_cluster_sb_BL_4_11, wire_in_cluster_sb_BL_3_11, wire_in_cluster_sb_BL_2_11, wire_in_cluster_sb_BL_1_11, wire_in_cluster_sb_BL_0_11 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_14, wire_in_cluster_sb_BL_14_14, wire_in_cluster_sb_BL_13_14, wire_in_cluster_sb_BL_12_14, wire_in_cluster_sb_BL_11_14, wire_in_cluster_sb_BL_10_14, wire_in_cluster_sb_BL_9_14, wire_in_cluster_sb_BL_8_14, wire_in_cluster_sb_BL_7_14, wire_in_cluster_sb_BL_6_14, wire_in_cluster_sb_BL_5_14, wire_in_cluster_sb_BL_4_14, wire_in_cluster_sb_BL_3_14, wire_in_cluster_sb_BL_2_14, wire_in_cluster_sb_BL_1_14, wire_in_cluster_sb_BL_0_14 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_14, wire_in_cluster_sb_BR_14_14, wire_in_cluster_sb_BR_13_14, wire_in_cluster_sb_BR_12_14, wire_in_cluster_sb_BR_11_14, wire_in_cluster_sb_BR_10_14, wire_in_cluster_sb_BR_9_14, wire_in_cluster_sb_BR_8_14, wire_in_cluster_sb_BR_7_14, wire_in_cluster_sb_BR_6_14, wire_in_cluster_sb_BR_5_14, wire_in_cluster_sb_BR_4_14, wire_in_cluster_sb_BR_3_14, wire_in_cluster_sb_BR_2_14, wire_in_cluster_sb_BR_1_14, wire_in_cluster_sb_BR_0_14 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_14, wire_in_cluster_sb_TL_14_14, wire_in_cluster_sb_TL_13_14, wire_in_cluster_sb_TL_12_14, wire_in_cluster_sb_TL_11_14, wire_in_cluster_sb_TL_10_14, wire_in_cluster_sb_TL_9_14, wire_in_cluster_sb_TL_8_14, wire_in_cluster_sb_TL_7_14, wire_in_cluster_sb_TL_6_14, wire_in_cluster_sb_TL_5_14, wire_in_cluster_sb_TL_4_14, wire_in_cluster_sb_TL_3_14, wire_in_cluster_sb_TL_2_14, wire_in_cluster_sb_TL_1_14, wire_in_cluster_sb_TL_0_14 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_15, wire_out_cluster_sb_TL_2_15, wire_out_cluster_sb_TL_1_15, wire_out_cluster_sb_TL_0_15 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_10, wire_out_cluster_sb_BR_2_10, wire_out_cluster_sb_BR_1_10, wire_out_cluster_sb_BR_0_10 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_11, wire_out_cluster_sb_BL_2_11, wire_out_cluster_sb_BL_1_11, wire_out_cluster_sb_BL_0_11 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_14, wire_out_cluster_sb_BL_2_14, wire_out_cluster_sb_BL_1_14, wire_out_cluster_sb_BL_0_14 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_14, wire_out_cluster_sb_BR_2_14, wire_out_cluster_sb_BR_1_14, wire_out_cluster_sb_BR_0_14 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_14, wire_out_cluster_sb_TL_2_14, wire_out_cluster_sb_TL_1_14, wire_out_cluster_sb_TL_0_14 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_18, wire_sb_bottom_input_10_18, wire_sb_bottom_input_9_18, wire_sb_bottom_input_8_18, wire_sb_bottom_input_7_18, wire_sb_bottom_input_6_18, wire_sb_bottom_input_5_18, wire_sb_bottom_input_4_18, wire_sb_bottom_input_3_18, wire_sb_bottom_input_2_18, wire_sb_bottom_input_1_18, wire_sb_bottom_input_0_18 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_18, wire_sb_bottom_output_10_18, wire_sb_bottom_output_9_18, wire_sb_bottom_output_8_18, wire_sb_bottom_output_7_18, wire_sb_bottom_output_6_18, wire_sb_bottom_output_5_18, wire_sb_bottom_output_4_18, wire_sb_bottom_output_3_18, wire_sb_bottom_output_2_18, wire_sb_bottom_output_1_18, wire_sb_bottom_output_0_18 } )
      , .sb_left_input( { wire_sb_left_input_11_14, wire_sb_left_input_10_14, wire_sb_left_input_9_14, wire_sb_left_input_8_14, wire_sb_left_input_7_14, wire_sb_left_input_6_14, wire_sb_left_input_5_14, wire_sb_left_input_4_14, wire_sb_left_input_3_14, wire_sb_left_input_2_14, wire_sb_left_input_1_14, wire_sb_left_input_0_14 } )
      , .sb_left_output( { wire_sb_left_output_11_14, wire_sb_left_output_10_14, wire_sb_left_output_9_14, wire_sb_left_output_8_14, wire_sb_left_output_7_14, wire_sb_left_output_6_14, wire_sb_left_output_5_14, wire_sb_left_output_4_14, wire_sb_left_output_3_14, wire_sb_left_output_2_14, wire_sb_left_output_1_14, wire_sb_left_output_0_14 } )
      , .sb_right_input( { wire_sb_left_output_11_15, wire_sb_left_output_10_15, wire_sb_left_output_9_15, wire_sb_left_output_8_15, wire_sb_left_output_7_15, wire_sb_left_output_6_15, wire_sb_left_output_5_15, wire_sb_left_output_4_15, wire_sb_left_output_3_15, wire_sb_left_output_2_15, wire_sb_left_output_1_15, wire_sb_left_output_0_15 } )
      , .sb_right_output( { wire_sb_left_input_11_15, wire_sb_left_input_10_15, wire_sb_left_input_9_15, wire_sb_left_input_8_15, wire_sb_left_input_7_15, wire_sb_left_input_6_15, wire_sb_left_input_5_15, wire_sb_left_input_4_15, wire_sb_left_input_3_15, wire_sb_left_input_2_15, wire_sb_left_input_1_15, wire_sb_left_input_0_15 } )
      , .sb_top_input( { wire_sb_bottom_output_11_13, wire_sb_bottom_output_10_13, wire_sb_bottom_output_9_13, wire_sb_bottom_output_8_13, wire_sb_bottom_output_7_13, wire_sb_bottom_output_6_13, wire_sb_bottom_output_5_13, wire_sb_bottom_output_4_13, wire_sb_bottom_output_3_13, wire_sb_bottom_output_2_13, wire_sb_bottom_output_1_13, wire_sb_bottom_output_0_13 } )
      , .sb_top_output( { wire_sb_bottom_input_11_13, wire_sb_bottom_input_10_13, wire_sb_bottom_input_9_13, wire_sb_bottom_input_8_13, wire_sb_bottom_input_7_13, wire_sb_bottom_input_6_13, wire_sb_bottom_input_5_13, wire_sb_bottom_input_4_13, wire_sb_bottom_input_3_13, wire_sb_bottom_input_2_13, wire_sb_bottom_input_1_13, wire_sb_bottom_input_0_13 } )
     );

TileInternal tile_I6(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[6] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_5, wire_in_cluster_sb_TL_14_5, wire_in_cluster_sb_TL_13_5, wire_in_cluster_sb_TL_12_5, wire_in_cluster_sb_TL_11_5, wire_in_cluster_sb_TL_10_5, wire_in_cluster_sb_TL_9_5, wire_in_cluster_sb_TL_8_5, wire_in_cluster_sb_TL_7_5, wire_in_cluster_sb_TL_6_5, wire_in_cluster_sb_TL_5_5, wire_in_cluster_sb_TL_4_5, wire_in_cluster_sb_TL_3_5, wire_in_cluster_sb_TL_2_5, wire_in_cluster_sb_TL_1_5, wire_in_cluster_sb_TL_0_5 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_0, wire_in_cluster_sb_BR_14_0, wire_in_cluster_sb_BR_13_0, wire_in_cluster_sb_BR_12_0, wire_in_cluster_sb_BR_11_0, wire_in_cluster_sb_BR_10_0, wire_in_cluster_sb_BR_9_0, wire_in_cluster_sb_BR_8_0, wire_in_cluster_sb_BR_7_0, wire_in_cluster_sb_BR_6_0, wire_in_cluster_sb_BR_5_0, wire_in_cluster_sb_BR_4_0, wire_in_cluster_sb_BR_3_0, wire_in_cluster_sb_BR_2_0, wire_in_cluster_sb_BR_1_0, wire_in_cluster_sb_BR_0_0 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_1, wire_in_cluster_sb_BL_14_1, wire_in_cluster_sb_BL_13_1, wire_in_cluster_sb_BL_12_1, wire_in_cluster_sb_BL_11_1, wire_in_cluster_sb_BL_10_1, wire_in_cluster_sb_BL_9_1, wire_in_cluster_sb_BL_8_1, wire_in_cluster_sb_BL_7_1, wire_in_cluster_sb_BL_6_1, wire_in_cluster_sb_BL_5_1, wire_in_cluster_sb_BL_4_1, wire_in_cluster_sb_BL_3_1, wire_in_cluster_sb_BL_2_1, wire_in_cluster_sb_BL_1_1, wire_in_cluster_sb_BL_0_1 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_4, wire_in_cluster_sb_BL_14_4, wire_in_cluster_sb_BL_13_4, wire_in_cluster_sb_BL_12_4, wire_in_cluster_sb_BL_11_4, wire_in_cluster_sb_BL_10_4, wire_in_cluster_sb_BL_9_4, wire_in_cluster_sb_BL_8_4, wire_in_cluster_sb_BL_7_4, wire_in_cluster_sb_BL_6_4, wire_in_cluster_sb_BL_5_4, wire_in_cluster_sb_BL_4_4, wire_in_cluster_sb_BL_3_4, wire_in_cluster_sb_BL_2_4, wire_in_cluster_sb_BL_1_4, wire_in_cluster_sb_BL_0_4 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_4, wire_in_cluster_sb_BR_14_4, wire_in_cluster_sb_BR_13_4, wire_in_cluster_sb_BR_12_4, wire_in_cluster_sb_BR_11_4, wire_in_cluster_sb_BR_10_4, wire_in_cluster_sb_BR_9_4, wire_in_cluster_sb_BR_8_4, wire_in_cluster_sb_BR_7_4, wire_in_cluster_sb_BR_6_4, wire_in_cluster_sb_BR_5_4, wire_in_cluster_sb_BR_4_4, wire_in_cluster_sb_BR_3_4, wire_in_cluster_sb_BR_2_4, wire_in_cluster_sb_BR_1_4, wire_in_cluster_sb_BR_0_4 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_4, wire_in_cluster_sb_TL_14_4, wire_in_cluster_sb_TL_13_4, wire_in_cluster_sb_TL_12_4, wire_in_cluster_sb_TL_11_4, wire_in_cluster_sb_TL_10_4, wire_in_cluster_sb_TL_9_4, wire_in_cluster_sb_TL_8_4, wire_in_cluster_sb_TL_7_4, wire_in_cluster_sb_TL_6_4, wire_in_cluster_sb_TL_5_4, wire_in_cluster_sb_TL_4_4, wire_in_cluster_sb_TL_3_4, wire_in_cluster_sb_TL_2_4, wire_in_cluster_sb_TL_1_4, wire_in_cluster_sb_TL_0_4 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_5, wire_out_cluster_sb_TL_2_5, wire_out_cluster_sb_TL_1_5, wire_out_cluster_sb_TL_0_5 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_0, wire_out_cluster_sb_BR_2_0, wire_out_cluster_sb_BR_1_0, wire_out_cluster_sb_BR_0_0 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_1, wire_out_cluster_sb_BL_2_1, wire_out_cluster_sb_BL_1_1, wire_out_cluster_sb_BL_0_1 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_4, wire_out_cluster_sb_BL_2_4, wire_out_cluster_sb_BL_1_4, wire_out_cluster_sb_BL_0_4 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_4, wire_out_cluster_sb_BR_2_4, wire_out_cluster_sb_BR_1_4, wire_out_cluster_sb_BR_0_4 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_4, wire_out_cluster_sb_TL_2_4, wire_out_cluster_sb_TL_1_4, wire_out_cluster_sb_TL_0_4 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_6, wire_sb_bottom_input_10_6, wire_sb_bottom_input_9_6, wire_sb_bottom_input_8_6, wire_sb_bottom_input_7_6, wire_sb_bottom_input_6_6, wire_sb_bottom_input_5_6, wire_sb_bottom_input_4_6, wire_sb_bottom_input_3_6, wire_sb_bottom_input_2_6, wire_sb_bottom_input_1_6, wire_sb_bottom_input_0_6 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_6, wire_sb_bottom_output_10_6, wire_sb_bottom_output_9_6, wire_sb_bottom_output_8_6, wire_sb_bottom_output_7_6, wire_sb_bottom_output_6_6, wire_sb_bottom_output_5_6, wire_sb_bottom_output_4_6, wire_sb_bottom_output_3_6, wire_sb_bottom_output_2_6, wire_sb_bottom_output_1_6, wire_sb_bottom_output_0_6 } )
      , .sb_left_input( { wire_sb_left_input_11_4, wire_sb_left_input_10_4, wire_sb_left_input_9_4, wire_sb_left_input_8_4, wire_sb_left_input_7_4, wire_sb_left_input_6_4, wire_sb_left_input_5_4, wire_sb_left_input_4_4, wire_sb_left_input_3_4, wire_sb_left_input_2_4, wire_sb_left_input_1_4, wire_sb_left_input_0_4 } )
      , .sb_left_output( { wire_sb_left_output_11_4, wire_sb_left_output_10_4, wire_sb_left_output_9_4, wire_sb_left_output_8_4, wire_sb_left_output_7_4, wire_sb_left_output_6_4, wire_sb_left_output_5_4, wire_sb_left_output_4_4, wire_sb_left_output_3_4, wire_sb_left_output_2_4, wire_sb_left_output_1_4, wire_sb_left_output_0_4 } )
      , .sb_right_input( { wire_sb_left_output_11_5, wire_sb_left_output_10_5, wire_sb_left_output_9_5, wire_sb_left_output_8_5, wire_sb_left_output_7_5, wire_sb_left_output_6_5, wire_sb_left_output_5_5, wire_sb_left_output_4_5, wire_sb_left_output_3_5, wire_sb_left_output_2_5, wire_sb_left_output_1_5, wire_sb_left_output_0_5 } )
      , .sb_right_output( { wire_sb_left_input_11_5, wire_sb_left_input_10_5, wire_sb_left_input_9_5, wire_sb_left_input_8_5, wire_sb_left_input_7_5, wire_sb_left_input_6_5, wire_sb_left_input_5_5, wire_sb_left_input_4_5, wire_sb_left_input_3_5, wire_sb_left_input_2_5, wire_sb_left_input_1_5, wire_sb_left_input_0_5 } )
      , .sb_top_input( { wire_sb_bottom_output_11_1, wire_sb_bottom_output_10_1, wire_sb_bottom_output_9_1, wire_sb_bottom_output_8_1, wire_sb_bottom_output_7_1, wire_sb_bottom_output_6_1, wire_sb_bottom_output_5_1, wire_sb_bottom_output_4_1, wire_sb_bottom_output_3_1, wire_sb_bottom_output_2_1, wire_sb_bottom_output_1_1, wire_sb_bottom_output_0_1 } )
      , .sb_top_output( { wire_sb_bottom_input_11_1, wire_sb_bottom_input_10_1, wire_sb_bottom_input_9_1, wire_sb_bottom_input_8_1, wire_sb_bottom_input_7_1, wire_sb_bottom_input_6_1, wire_sb_bottom_input_5_1, wire_sb_bottom_input_4_1, wire_sb_bottom_input_3_1, wire_sb_bottom_input_2_1, wire_sb_bottom_input_1_1, wire_sb_bottom_input_0_1 } )
     );

TileInternal tile_I7(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[7] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_6, wire_in_cluster_sb_TL_14_6, wire_in_cluster_sb_TL_13_6, wire_in_cluster_sb_TL_12_6, wire_in_cluster_sb_TL_11_6, wire_in_cluster_sb_TL_10_6, wire_in_cluster_sb_TL_9_6, wire_in_cluster_sb_TL_8_6, wire_in_cluster_sb_TL_7_6, wire_in_cluster_sb_TL_6_6, wire_in_cluster_sb_TL_5_6, wire_in_cluster_sb_TL_4_6, wire_in_cluster_sb_TL_3_6, wire_in_cluster_sb_TL_2_6, wire_in_cluster_sb_TL_1_6, wire_in_cluster_sb_TL_0_6 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_1, wire_in_cluster_sb_BR_14_1, wire_in_cluster_sb_BR_13_1, wire_in_cluster_sb_BR_12_1, wire_in_cluster_sb_BR_11_1, wire_in_cluster_sb_BR_10_1, wire_in_cluster_sb_BR_9_1, wire_in_cluster_sb_BR_8_1, wire_in_cluster_sb_BR_7_1, wire_in_cluster_sb_BR_6_1, wire_in_cluster_sb_BR_5_1, wire_in_cluster_sb_BR_4_1, wire_in_cluster_sb_BR_3_1, wire_in_cluster_sb_BR_2_1, wire_in_cluster_sb_BR_1_1, wire_in_cluster_sb_BR_0_1 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_2, wire_in_cluster_sb_BL_14_2, wire_in_cluster_sb_BL_13_2, wire_in_cluster_sb_BL_12_2, wire_in_cluster_sb_BL_11_2, wire_in_cluster_sb_BL_10_2, wire_in_cluster_sb_BL_9_2, wire_in_cluster_sb_BL_8_2, wire_in_cluster_sb_BL_7_2, wire_in_cluster_sb_BL_6_2, wire_in_cluster_sb_BL_5_2, wire_in_cluster_sb_BL_4_2, wire_in_cluster_sb_BL_3_2, wire_in_cluster_sb_BL_2_2, wire_in_cluster_sb_BL_1_2, wire_in_cluster_sb_BL_0_2 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_5, wire_in_cluster_sb_BL_14_5, wire_in_cluster_sb_BL_13_5, wire_in_cluster_sb_BL_12_5, wire_in_cluster_sb_BL_11_5, wire_in_cluster_sb_BL_10_5, wire_in_cluster_sb_BL_9_5, wire_in_cluster_sb_BL_8_5, wire_in_cluster_sb_BL_7_5, wire_in_cluster_sb_BL_6_5, wire_in_cluster_sb_BL_5_5, wire_in_cluster_sb_BL_4_5, wire_in_cluster_sb_BL_3_5, wire_in_cluster_sb_BL_2_5, wire_in_cluster_sb_BL_1_5, wire_in_cluster_sb_BL_0_5 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_5, wire_in_cluster_sb_BR_14_5, wire_in_cluster_sb_BR_13_5, wire_in_cluster_sb_BR_12_5, wire_in_cluster_sb_BR_11_5, wire_in_cluster_sb_BR_10_5, wire_in_cluster_sb_BR_9_5, wire_in_cluster_sb_BR_8_5, wire_in_cluster_sb_BR_7_5, wire_in_cluster_sb_BR_6_5, wire_in_cluster_sb_BR_5_5, wire_in_cluster_sb_BR_4_5, wire_in_cluster_sb_BR_3_5, wire_in_cluster_sb_BR_2_5, wire_in_cluster_sb_BR_1_5, wire_in_cluster_sb_BR_0_5 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_5, wire_in_cluster_sb_TL_14_5, wire_in_cluster_sb_TL_13_5, wire_in_cluster_sb_TL_12_5, wire_in_cluster_sb_TL_11_5, wire_in_cluster_sb_TL_10_5, wire_in_cluster_sb_TL_9_5, wire_in_cluster_sb_TL_8_5, wire_in_cluster_sb_TL_7_5, wire_in_cluster_sb_TL_6_5, wire_in_cluster_sb_TL_5_5, wire_in_cluster_sb_TL_4_5, wire_in_cluster_sb_TL_3_5, wire_in_cluster_sb_TL_2_5, wire_in_cluster_sb_TL_1_5, wire_in_cluster_sb_TL_0_5 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_6, wire_out_cluster_sb_TL_2_6, wire_out_cluster_sb_TL_1_6, wire_out_cluster_sb_TL_0_6 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_1, wire_out_cluster_sb_BR_2_1, wire_out_cluster_sb_BR_1_1, wire_out_cluster_sb_BR_0_1 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_2, wire_out_cluster_sb_BL_2_2, wire_out_cluster_sb_BL_1_2, wire_out_cluster_sb_BL_0_2 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_5, wire_out_cluster_sb_BL_2_5, wire_out_cluster_sb_BL_1_5, wire_out_cluster_sb_BL_0_5 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_5, wire_out_cluster_sb_BR_2_5, wire_out_cluster_sb_BR_1_5, wire_out_cluster_sb_BR_0_5 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_5, wire_out_cluster_sb_TL_2_5, wire_out_cluster_sb_TL_1_5, wire_out_cluster_sb_TL_0_5 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_7, wire_sb_bottom_input_10_7, wire_sb_bottom_input_9_7, wire_sb_bottom_input_8_7, wire_sb_bottom_input_7_7, wire_sb_bottom_input_6_7, wire_sb_bottom_input_5_7, wire_sb_bottom_input_4_7, wire_sb_bottom_input_3_7, wire_sb_bottom_input_2_7, wire_sb_bottom_input_1_7, wire_sb_bottom_input_0_7 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_7, wire_sb_bottom_output_10_7, wire_sb_bottom_output_9_7, wire_sb_bottom_output_8_7, wire_sb_bottom_output_7_7, wire_sb_bottom_output_6_7, wire_sb_bottom_output_5_7, wire_sb_bottom_output_4_7, wire_sb_bottom_output_3_7, wire_sb_bottom_output_2_7, wire_sb_bottom_output_1_7, wire_sb_bottom_output_0_7 } )
      , .sb_left_input( { wire_sb_left_input_11_5, wire_sb_left_input_10_5, wire_sb_left_input_9_5, wire_sb_left_input_8_5, wire_sb_left_input_7_5, wire_sb_left_input_6_5, wire_sb_left_input_5_5, wire_sb_left_input_4_5, wire_sb_left_input_3_5, wire_sb_left_input_2_5, wire_sb_left_input_1_5, wire_sb_left_input_0_5 } )
      , .sb_left_output( { wire_sb_left_output_11_5, wire_sb_left_output_10_5, wire_sb_left_output_9_5, wire_sb_left_output_8_5, wire_sb_left_output_7_5, wire_sb_left_output_6_5, wire_sb_left_output_5_5, wire_sb_left_output_4_5, wire_sb_left_output_3_5, wire_sb_left_output_2_5, wire_sb_left_output_1_5, wire_sb_left_output_0_5 } )
      , .sb_right_input( { wire_sb_left_output_11_6, wire_sb_left_output_10_6, wire_sb_left_output_9_6, wire_sb_left_output_8_6, wire_sb_left_output_7_6, wire_sb_left_output_6_6, wire_sb_left_output_5_6, wire_sb_left_output_4_6, wire_sb_left_output_3_6, wire_sb_left_output_2_6, wire_sb_left_output_1_6, wire_sb_left_output_0_6 } )
      , .sb_right_output( { wire_sb_left_input_11_6, wire_sb_left_input_10_6, wire_sb_left_input_9_6, wire_sb_left_input_8_6, wire_sb_left_input_7_6, wire_sb_left_input_6_6, wire_sb_left_input_5_6, wire_sb_left_input_4_6, wire_sb_left_input_3_6, wire_sb_left_input_2_6, wire_sb_left_input_1_6, wire_sb_left_input_0_6 } )
      , .sb_top_input( { wire_sb_bottom_output_11_2, wire_sb_bottom_output_10_2, wire_sb_bottom_output_9_2, wire_sb_bottom_output_8_2, wire_sb_bottom_output_7_2, wire_sb_bottom_output_6_2, wire_sb_bottom_output_5_2, wire_sb_bottom_output_4_2, wire_sb_bottom_output_3_2, wire_sb_bottom_output_2_2, wire_sb_bottom_output_1_2, wire_sb_bottom_output_0_2 } )
      , .sb_top_output( { wire_sb_bottom_input_11_2, wire_sb_bottom_input_10_2, wire_sb_bottom_input_9_2, wire_sb_bottom_input_8_2, wire_sb_bottom_input_7_2, wire_sb_bottom_input_6_2, wire_sb_bottom_input_5_2, wire_sb_bottom_input_4_2, wire_sb_bottom_input_3_2, wire_sb_bottom_input_2_2, wire_sb_bottom_input_1_2, wire_sb_bottom_input_0_2 } )
     );

TileInternal tile_I8(
        .clock( clock )
      , .conf( conf )
      , .reset( reset )
      , .select_tile( w_SELECT_TILE_0[8] )
      , .address_tile( { w_ADDRESS_TILE_0[9], w_ADDRESS_TILE_0[8], w_ADDRESS_TILE_0[7], w_ADDRESS_TILE_0[6], w_ADDRESS_TILE_0[5], w_ADDRESS_TILE_0[4], w_ADDRESS_TILE_0[3], w_ADDRESS_TILE_0[2], w_ADDRESS_TILE_0[1], w_ADDRESS_TILE_0[0] } )
      , .data_tile( { data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0] } )
      , .in_cluster_BR( { wire_in_cluster_sb_TL_15_7, wire_in_cluster_sb_TL_14_7, wire_in_cluster_sb_TL_13_7, wire_in_cluster_sb_TL_12_7, wire_in_cluster_sb_TL_11_7, wire_in_cluster_sb_TL_10_7, wire_in_cluster_sb_TL_9_7, wire_in_cluster_sb_TL_8_7, wire_in_cluster_sb_TL_7_7, wire_in_cluster_sb_TL_6_7, wire_in_cluster_sb_TL_5_7, wire_in_cluster_sb_TL_4_7, wire_in_cluster_sb_TL_3_7, wire_in_cluster_sb_TL_2_7, wire_in_cluster_sb_TL_1_7, wire_in_cluster_sb_TL_0_7 } )
      , .in_cluster_TL( { wire_in_cluster_sb_BR_15_2, wire_in_cluster_sb_BR_14_2, wire_in_cluster_sb_BR_13_2, wire_in_cluster_sb_BR_12_2, wire_in_cluster_sb_BR_11_2, wire_in_cluster_sb_BR_10_2, wire_in_cluster_sb_BR_9_2, wire_in_cluster_sb_BR_8_2, wire_in_cluster_sb_BR_7_2, wire_in_cluster_sb_BR_6_2, wire_in_cluster_sb_BR_5_2, wire_in_cluster_sb_BR_4_2, wire_in_cluster_sb_BR_3_2, wire_in_cluster_sb_BR_2_2, wire_in_cluster_sb_BR_1_2, wire_in_cluster_sb_BR_0_2 } )
      , .in_cluster_TR( { wire_in_cluster_sb_BL_15_3, wire_in_cluster_sb_BL_14_3, wire_in_cluster_sb_BL_13_3, wire_in_cluster_sb_BL_12_3, wire_in_cluster_sb_BL_11_3, wire_in_cluster_sb_BL_10_3, wire_in_cluster_sb_BL_9_3, wire_in_cluster_sb_BL_8_3, wire_in_cluster_sb_BL_7_3, wire_in_cluster_sb_BL_6_3, wire_in_cluster_sb_BL_5_3, wire_in_cluster_sb_BL_4_3, wire_in_cluster_sb_BL_3_3, wire_in_cluster_sb_BL_2_3, wire_in_cluster_sb_BL_1_3, wire_in_cluster_sb_BL_0_3 } )
      , .in_cluster_sb_BL( { wire_in_cluster_sb_BL_15_6, wire_in_cluster_sb_BL_14_6, wire_in_cluster_sb_BL_13_6, wire_in_cluster_sb_BL_12_6, wire_in_cluster_sb_BL_11_6, wire_in_cluster_sb_BL_10_6, wire_in_cluster_sb_BL_9_6, wire_in_cluster_sb_BL_8_6, wire_in_cluster_sb_BL_7_6, wire_in_cluster_sb_BL_6_6, wire_in_cluster_sb_BL_5_6, wire_in_cluster_sb_BL_4_6, wire_in_cluster_sb_BL_3_6, wire_in_cluster_sb_BL_2_6, wire_in_cluster_sb_BL_1_6, wire_in_cluster_sb_BL_0_6 } )
      , .in_cluster_sb_BR( { wire_in_cluster_sb_BR_15_6, wire_in_cluster_sb_BR_14_6, wire_in_cluster_sb_BR_13_6, wire_in_cluster_sb_BR_12_6, wire_in_cluster_sb_BR_11_6, wire_in_cluster_sb_BR_10_6, wire_in_cluster_sb_BR_9_6, wire_in_cluster_sb_BR_8_6, wire_in_cluster_sb_BR_7_6, wire_in_cluster_sb_BR_6_6, wire_in_cluster_sb_BR_5_6, wire_in_cluster_sb_BR_4_6, wire_in_cluster_sb_BR_3_6, wire_in_cluster_sb_BR_2_6, wire_in_cluster_sb_BR_1_6, wire_in_cluster_sb_BR_0_6 } )
      , .in_cluster_sb_TL( { wire_in_cluster_sb_TL_15_6, wire_in_cluster_sb_TL_14_6, wire_in_cluster_sb_TL_13_6, wire_in_cluster_sb_TL_12_6, wire_in_cluster_sb_TL_11_6, wire_in_cluster_sb_TL_10_6, wire_in_cluster_sb_TL_9_6, wire_in_cluster_sb_TL_8_6, wire_in_cluster_sb_TL_7_6, wire_in_cluster_sb_TL_6_6, wire_in_cluster_sb_TL_5_6, wire_in_cluster_sb_TL_4_6, wire_in_cluster_sb_TL_3_6, wire_in_cluster_sb_TL_2_6, wire_in_cluster_sb_TL_1_6, wire_in_cluster_sb_TL_0_6 } )
      , .out_cluster_BR( { wire_out_cluster_sb_TL_3_7, wire_out_cluster_sb_TL_2_7, wire_out_cluster_sb_TL_1_7, wire_out_cluster_sb_TL_0_7 } )
      , .out_cluster_TL( { wire_out_cluster_sb_BR_3_2, wire_out_cluster_sb_BR_2_2, wire_out_cluster_sb_BR_1_2, wire_out_cluster_sb_BR_0_2 } )
      , .out_cluster_TR( { wire_out_cluster_sb_BL_3_3, wire_out_cluster_sb_BL_2_3, wire_out_cluster_sb_BL_1_3, wire_out_cluster_sb_BL_0_3 } )
      , .out_cluster_sb_BL( { wire_out_cluster_sb_BL_3_6, wire_out_cluster_sb_BL_2_6, wire_out_cluster_sb_BL_1_6, wire_out_cluster_sb_BL_0_6 } )
      , .out_cluster_sb_BR( { wire_out_cluster_sb_BR_3_6, wire_out_cluster_sb_BR_2_6, wire_out_cluster_sb_BR_1_6, wire_out_cluster_sb_BR_0_6 } )
      , .out_cluster_sb_TL( { wire_out_cluster_sb_TL_3_6, wire_out_cluster_sb_TL_2_6, wire_out_cluster_sb_TL_1_6, wire_out_cluster_sb_TL_0_6 } )
      , .sb_bottom_input( { wire_sb_bottom_input_11_8, wire_sb_bottom_input_10_8, wire_sb_bottom_input_9_8, wire_sb_bottom_input_8_8, wire_sb_bottom_input_7_8, wire_sb_bottom_input_6_8, wire_sb_bottom_input_5_8, wire_sb_bottom_input_4_8, wire_sb_bottom_input_3_8, wire_sb_bottom_input_2_8, wire_sb_bottom_input_1_8, wire_sb_bottom_input_0_8 } )
      , .sb_bottom_output( { wire_sb_bottom_output_11_8, wire_sb_bottom_output_10_8, wire_sb_bottom_output_9_8, wire_sb_bottom_output_8_8, wire_sb_bottom_output_7_8, wire_sb_bottom_output_6_8, wire_sb_bottom_output_5_8, wire_sb_bottom_output_4_8, wire_sb_bottom_output_3_8, wire_sb_bottom_output_2_8, wire_sb_bottom_output_1_8, wire_sb_bottom_output_0_8 } )
      , .sb_left_input( { wire_sb_left_input_11_6, wire_sb_left_input_10_6, wire_sb_left_input_9_6, wire_sb_left_input_8_6, wire_sb_left_input_7_6, wire_sb_left_input_6_6, wire_sb_left_input_5_6, wire_sb_left_input_4_6, wire_sb_left_input_3_6, wire_sb_left_input_2_6, wire_sb_left_input_1_6, wire_sb_left_input_0_6 } )
      , .sb_left_output( { wire_sb_left_output_11_6, wire_sb_left_output_10_6, wire_sb_left_output_9_6, wire_sb_left_output_8_6, wire_sb_left_output_7_6, wire_sb_left_output_6_6, wire_sb_left_output_5_6, wire_sb_left_output_4_6, wire_sb_left_output_3_6, wire_sb_left_output_2_6, wire_sb_left_output_1_6, wire_sb_left_output_0_6 } )
      , .sb_right_input( { wire_sb_left_output_11_7, wire_sb_left_output_10_7, wire_sb_left_output_9_7, wire_sb_left_output_8_7, wire_sb_left_output_7_7, wire_sb_left_output_6_7, wire_sb_left_output_5_7, wire_sb_left_output_4_7, wire_sb_left_output_3_7, wire_sb_left_output_2_7, wire_sb_left_output_1_7, wire_sb_left_output_0_7 } )
      , .sb_right_output( { wire_sb_left_input_11_7, wire_sb_left_input_10_7, wire_sb_left_input_9_7, wire_sb_left_input_8_7, wire_sb_left_input_7_7, wire_sb_left_input_6_7, wire_sb_left_input_5_7, wire_sb_left_input_4_7, wire_sb_left_input_3_7, wire_sb_left_input_2_7, wire_sb_left_input_1_7, wire_sb_left_input_0_7 } )
      , .sb_top_input( { wire_sb_bottom_output_11_3, wire_sb_bottom_output_10_3, wire_sb_bottom_output_9_3, wire_sb_bottom_output_8_3, wire_sb_bottom_output_7_3, wire_sb_bottom_output_6_3, wire_sb_bottom_output_5_3, wire_sb_bottom_output_4_3, wire_sb_bottom_output_3_3, wire_sb_bottom_output_2_3, wire_sb_bottom_output_1_3, wire_sb_bottom_output_0_3 } )
      , .sb_top_output( { wire_sb_bottom_input_11_3, wire_sb_bottom_input_10_3, wire_sb_bottom_input_9_3, wire_sb_bottom_input_8_3, wire_sb_bottom_input_7_3, wire_sb_bottom_input_6_3, wire_sb_bottom_input_5_3, wire_sb_bottom_input_4_3, wire_sb_bottom_input_3_3, wire_sb_bottom_input_2_3, wire_sb_bottom_input_1_3, wire_sb_bottom_input_0_3 } )
     );


endmodule
