`timescale 1 ns/1 ps

module cluster_1(
     func_ck1
   , conf_ck1
   , selector1
   , reset1
   , input_tree1
   , output_tree1
   , cluster_data1
   , address1
  );


input   func_ck1;
wire func_ck1;
input   conf_ck1;
wire conf_ck1;
input   selector1;
wire selector1;
input   reset1;
wire reset1;
input   [63:0] input_tree1;
wire [63:0] input_tree1;
output  [15:0] output_tree1;
wire [15:0] output_tree1;
input   [7:0] cluster_data1;
wire [7:0] cluster_data1;
input   [8:0] address1;
wire [8:0] address1;

wire wire_INPUTS_0_0;
wire wire_INPUTS_0_1;
wire wire_INPUTS_0_10;
wire wire_INPUTS_0_11;
wire wire_INPUTS_0_12;
wire wire_INPUTS_0_13;
wire wire_INPUTS_0_14;
wire wire_INPUTS_0_15;
wire wire_INPUTS_0_2;
wire wire_INPUTS_0_3;
wire wire_INPUTS_0_4;
wire wire_INPUTS_0_5;
wire wire_INPUTS_0_6;
wire wire_INPUTS_0_7;
wire wire_INPUTS_0_8;
wire wire_INPUTS_0_9;
wire [5:0] w_ADDRESS_LEVEL_D_0;
wire [3:0] w_SELECT_LEVEL_D_0;
wire [63:0] w_STROBE_DMSB_0;
wire [31:0] w_STROBE_UMSB_0;
wire [3:0] w_dmsb0_OUTPUTS;
wire [3:0] w_dmsb10_OUTPUTS;
wire [3:0] w_dmsb11_OUTPUTS;
wire [3:0] w_dmsb12_OUTPUTS;
wire [3:0] w_dmsb13_OUTPUTS;
wire [3:0] w_dmsb14_OUTPUTS;
wire [3:0] w_dmsb15_OUTPUTS;
wire [3:0] w_dmsb1_OUTPUTS;
wire [3:0] w_dmsb2_OUTPUTS;
wire [3:0] w_dmsb3_OUTPUTS;
wire [3:0] w_dmsb4_OUTPUTS;
wire [3:0] w_dmsb5_OUTPUTS;
wire [3:0] w_dmsb6_OUTPUTS;
wire [3:0] w_dmsb7_OUTPUTS;
wire [3:0] w_dmsb8_OUTPUTS;
wire [3:0] w_dmsb9_OUTPUTS;
wire [3:0] w_umsb0_INPUTS;
wire [3:0] w_umsb1_INPUTS;
wire [3:0] w_umsb2_INPUTS;
wire [3:0] w_umsb3_INPUTS;

cluster_0 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop(
        .conf_ck0( conf_ck1 )
      , .func_ck0( func_ck1 )
      , .reset0( reset1 )
      , .selector0( w_SELECT_LEVEL_D_0[0] )
      , .address0( { address1[5], address1[4], address1[3], address1[2], address1[1], address1[0] } )
      , .cluster_data0( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .cluster_inputs0( { w_dmsb15_OUTPUTS[0], w_dmsb11_OUTPUTS[0], w_dmsb7_OUTPUTS[0], w_dmsb3_OUTPUTS[0], w_dmsb14_OUTPUTS[0], w_dmsb10_OUTPUTS[0], w_dmsb6_OUTPUTS[0], w_dmsb2_OUTPUTS[0], w_dmsb13_OUTPUTS[0], w_dmsb9_OUTPUTS[0], w_dmsb5_OUTPUTS[0], w_dmsb1_OUTPUTS[0], w_dmsb12_OUTPUTS[0], w_dmsb8_OUTPUTS[0], w_dmsb4_OUTPUTS[0], w_dmsb0_OUTPUTS[0] } )
      , .cluster_outputs0( { w_umsb3_INPUTS[0], w_umsb2_INPUTS[0], w_umsb1_INPUTS[0], w_umsb0_INPUTS[0] } )
      , .input_tree0( { input_tree1[15], input_tree1[14], input_tree1[13], input_tree1[12], input_tree1[11], input_tree1[10], input_tree1[9], input_tree1[8], input_tree1[7], input_tree1[6], input_tree1[5], input_tree1[4], input_tree1[3], input_tree1[2], input_tree1[1], input_tree1[0] } )
      , .output_tree0( { output_tree1[3], output_tree1[2], output_tree1[1], output_tree1[0] } )
     );

cluster_0 cluster_0_instance_cluster1_TileBoundaryTop_TileBoundaryTop(
        .conf_ck0( conf_ck1 )
      , .func_ck0( func_ck1 )
      , .reset0( reset1 )
      , .selector0( w_SELECT_LEVEL_D_0[1] )
      , .address0( { address1[5], address1[4], address1[3], address1[2], address1[1], address1[0] } )
      , .cluster_data0( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .cluster_inputs0( { w_dmsb15_OUTPUTS[1], w_dmsb11_OUTPUTS[1], w_dmsb7_OUTPUTS[1], w_dmsb3_OUTPUTS[1], w_dmsb14_OUTPUTS[1], w_dmsb10_OUTPUTS[1], w_dmsb6_OUTPUTS[1], w_dmsb2_OUTPUTS[1], w_dmsb13_OUTPUTS[1], w_dmsb9_OUTPUTS[1], w_dmsb5_OUTPUTS[1], w_dmsb1_OUTPUTS[1], w_dmsb12_OUTPUTS[1], w_dmsb8_OUTPUTS[1], w_dmsb4_OUTPUTS[1], w_dmsb0_OUTPUTS[1] } )
      , .cluster_outputs0( { w_umsb3_INPUTS[1], w_umsb2_INPUTS[1], w_umsb1_INPUTS[1], w_umsb0_INPUTS[1] } )
      , .input_tree0( { input_tree1[31], input_tree1[30], input_tree1[29], input_tree1[28], input_tree1[27], input_tree1[26], input_tree1[25], input_tree1[24], input_tree1[23], input_tree1[22], input_tree1[21], input_tree1[20], input_tree1[19], input_tree1[18], input_tree1[17], input_tree1[16] } )
      , .output_tree0( { output_tree1[7], output_tree1[6], output_tree1[5], output_tree1[4] } )
     );

cluster_0 cluster_0_instance_cluster2_TileBoundaryTop_TileBoundaryTop(
        .conf_ck0( conf_ck1 )
      , .func_ck0( func_ck1 )
      , .reset0( reset1 )
      , .selector0( w_SELECT_LEVEL_D_0[2] )
      , .address0( { address1[5], address1[4], address1[3], address1[2], address1[1], address1[0] } )
      , .cluster_data0( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .cluster_inputs0( { w_dmsb15_OUTPUTS[2], w_dmsb11_OUTPUTS[2], w_dmsb7_OUTPUTS[2], w_dmsb3_OUTPUTS[2], w_dmsb14_OUTPUTS[2], w_dmsb10_OUTPUTS[2], w_dmsb6_OUTPUTS[2], w_dmsb2_OUTPUTS[2], w_dmsb13_OUTPUTS[2], w_dmsb9_OUTPUTS[2], w_dmsb5_OUTPUTS[2], w_dmsb1_OUTPUTS[2], w_dmsb12_OUTPUTS[2], w_dmsb8_OUTPUTS[2], w_dmsb4_OUTPUTS[2], w_dmsb0_OUTPUTS[2] } )
      , .cluster_outputs0( { w_umsb3_INPUTS[2], w_umsb2_INPUTS[2], w_umsb1_INPUTS[2], w_umsb0_INPUTS[2] } )
      , .input_tree0( { input_tree1[47], input_tree1[46], input_tree1[45], input_tree1[44], input_tree1[43], input_tree1[42], input_tree1[41], input_tree1[40], input_tree1[39], input_tree1[38], input_tree1[37], input_tree1[36], input_tree1[35], input_tree1[34], input_tree1[33], input_tree1[32] } )
      , .output_tree0( { output_tree1[11], output_tree1[10], output_tree1[9], output_tree1[8] } )
     );

cluster_0 cluster_0_instance_cluster3_TileBoundaryTop_TileBoundaryTop(
        .conf_ck0( conf_ck1 )
      , .func_ck0( func_ck1 )
      , .reset0( reset1 )
      , .selector0( w_SELECT_LEVEL_D_0[3] )
      , .address0( { address1[5], address1[4], address1[3], address1[2], address1[1], address1[0] } )
      , .cluster_data0( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .cluster_inputs0( { w_dmsb15_OUTPUTS[3], w_dmsb11_OUTPUTS[3], w_dmsb7_OUTPUTS[3], w_dmsb3_OUTPUTS[3], w_dmsb14_OUTPUTS[3], w_dmsb10_OUTPUTS[3], w_dmsb6_OUTPUTS[3], w_dmsb2_OUTPUTS[3], w_dmsb13_OUTPUTS[3], w_dmsb9_OUTPUTS[3], w_dmsb5_OUTPUTS[3], w_dmsb1_OUTPUTS[3], w_dmsb12_OUTPUTS[3], w_dmsb8_OUTPUTS[3], w_dmsb4_OUTPUTS[3], w_dmsb0_OUTPUTS[3] } )
      , .cluster_outputs0( { w_umsb3_INPUTS[3], w_umsb2_INPUTS[3], w_umsb1_INPUTS[3], w_umsb0_INPUTS[3] } )
      , .input_tree0( { input_tree1[63], input_tree1[62], input_tree1[61], input_tree1[60], input_tree1[59], input_tree1[58], input_tree1[57], input_tree1[56], input_tree1[55], input_tree1[54], input_tree1[53], input_tree1[52], input_tree1[51], input_tree1[50], input_tree1[49], input_tree1[48] } )
      , .output_tree0( { output_tree1[15], output_tree1[14], output_tree1[13], output_tree1[12] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_0(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_0 } )
      , .OUTPUTS( { w_dmsb0_OUTPUTS[3], w_dmsb0_OUTPUTS[2], w_dmsb0_OUTPUTS[1], w_dmsb0_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[3], w_STROBE_DMSB_0[2], w_STROBE_DMSB_0[1], w_STROBE_DMSB_0[0] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_1(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_1 } )
      , .OUTPUTS( { w_dmsb1_OUTPUTS[3], w_dmsb1_OUTPUTS[2], w_dmsb1_OUTPUTS[1], w_dmsb1_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[7], w_STROBE_DMSB_0[6], w_STROBE_DMSB_0[5], w_STROBE_DMSB_0[4] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_10(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_10 } )
      , .OUTPUTS( { w_dmsb10_OUTPUTS[3], w_dmsb10_OUTPUTS[2], w_dmsb10_OUTPUTS[1], w_dmsb10_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[43], w_STROBE_DMSB_0[42], w_STROBE_DMSB_0[41], w_STROBE_DMSB_0[40] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_11(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_11 } )
      , .OUTPUTS( { w_dmsb11_OUTPUTS[3], w_dmsb11_OUTPUTS[2], w_dmsb11_OUTPUTS[1], w_dmsb11_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[47], w_STROBE_DMSB_0[46], w_STROBE_DMSB_0[45], w_STROBE_DMSB_0[44] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_12(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_12 } )
      , .OUTPUTS( { w_dmsb12_OUTPUTS[3], w_dmsb12_OUTPUTS[2], w_dmsb12_OUTPUTS[1], w_dmsb12_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[51], w_STROBE_DMSB_0[50], w_STROBE_DMSB_0[49], w_STROBE_DMSB_0[48] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_13(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_13 } )
      , .OUTPUTS( { w_dmsb13_OUTPUTS[3], w_dmsb13_OUTPUTS[2], w_dmsb13_OUTPUTS[1], w_dmsb13_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[55], w_STROBE_DMSB_0[54], w_STROBE_DMSB_0[53], w_STROBE_DMSB_0[52] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_14(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_14 } )
      , .OUTPUTS( { w_dmsb14_OUTPUTS[3], w_dmsb14_OUTPUTS[2], w_dmsb14_OUTPUTS[1], w_dmsb14_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[59], w_STROBE_DMSB_0[58], w_STROBE_DMSB_0[57], w_STROBE_DMSB_0[56] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_15(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_15 } )
      , .OUTPUTS( { w_dmsb15_OUTPUTS[3], w_dmsb15_OUTPUTS[2], w_dmsb15_OUTPUTS[1], w_dmsb15_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[63], w_STROBE_DMSB_0[62], w_STROBE_DMSB_0[61], w_STROBE_DMSB_0[60] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_2(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_2 } )
      , .OUTPUTS( { w_dmsb2_OUTPUTS[3], w_dmsb2_OUTPUTS[2], w_dmsb2_OUTPUTS[1], w_dmsb2_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[11], w_STROBE_DMSB_0[10], w_STROBE_DMSB_0[9], w_STROBE_DMSB_0[8] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_3(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_3 } )
      , .OUTPUTS( { w_dmsb3_OUTPUTS[3], w_dmsb3_OUTPUTS[2], w_dmsb3_OUTPUTS[1], w_dmsb3_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[15], w_STROBE_DMSB_0[14], w_STROBE_DMSB_0[13], w_STROBE_DMSB_0[12] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_4(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_4 } )
      , .OUTPUTS( { w_dmsb4_OUTPUTS[3], w_dmsb4_OUTPUTS[2], w_dmsb4_OUTPUTS[1], w_dmsb4_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[19], w_STROBE_DMSB_0[18], w_STROBE_DMSB_0[17], w_STROBE_DMSB_0[16] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_5(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_5 } )
      , .OUTPUTS( { w_dmsb5_OUTPUTS[3], w_dmsb5_OUTPUTS[2], w_dmsb5_OUTPUTS[1], w_dmsb5_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[23], w_STROBE_DMSB_0[22], w_STROBE_DMSB_0[21], w_STROBE_DMSB_0[20] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_6(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_6 } )
      , .OUTPUTS( { w_dmsb6_OUTPUTS[3], w_dmsb6_OUTPUTS[2], w_dmsb6_OUTPUTS[1], w_dmsb6_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[27], w_STROBE_DMSB_0[26], w_STROBE_DMSB_0[25], w_STROBE_DMSB_0[24] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_7(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_7 } )
      , .OUTPUTS( { w_dmsb7_OUTPUTS[3], w_dmsb7_OUTPUTS[2], w_dmsb7_OUTPUTS[1], w_dmsb7_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[31], w_STROBE_DMSB_0[30], w_STROBE_DMSB_0[29], w_STROBE_DMSB_0[28] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_8(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_8 } )
      , .OUTPUTS( { w_dmsb8_OUTPUTS[3], w_dmsb8_OUTPUTS[2], w_dmsb8_OUTPUTS[1], w_dmsb8_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[35], w_STROBE_DMSB_0[34], w_STROBE_DMSB_0[33], w_STROBE_DMSB_0[32] } )
     );

DMSB_NB_INPUTS_1_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_4 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_dmsb_9(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { wire_INPUTS_0_9 } )
      , .OUTPUTS( { w_dmsb9_OUTPUTS[3], w_dmsb9_OUTPUTS[2], w_dmsb9_OUTPUTS[1], w_dmsb9_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[39], w_STROBE_DMSB_0[38], w_STROBE_DMSB_0[37], w_STROBE_DMSB_0[36] } )
     );

UMSB_NB_INPUTS_4_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_8 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_umsb_0(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { w_umsb0_INPUTS[3], w_umsb0_INPUTS[2], w_umsb0_INPUTS[1], w_umsb0_INPUTS[0] } )
      , .OUTPUTS( { wire_INPUTS_0_3, wire_INPUTS_0_2, wire_INPUTS_0_1, wire_INPUTS_0_0 } )
      , .STROBE( { w_STROBE_UMSB_0[7], w_STROBE_UMSB_0[6], w_STROBE_UMSB_0[5], w_STROBE_UMSB_0[4], w_STROBE_UMSB_0[3], w_STROBE_UMSB_0[2], w_STROBE_UMSB_0[1], w_STROBE_UMSB_0[0] } )
     );

UMSB_NB_INPUTS_4_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_8 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_umsb_1(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { w_umsb1_INPUTS[3], w_umsb1_INPUTS[2], w_umsb1_INPUTS[1], w_umsb1_INPUTS[0] } )
      , .OUTPUTS( { wire_INPUTS_0_7, wire_INPUTS_0_6, wire_INPUTS_0_5, wire_INPUTS_0_4 } )
      , .STROBE( { w_STROBE_UMSB_0[15], w_STROBE_UMSB_0[14], w_STROBE_UMSB_0[13], w_STROBE_UMSB_0[12], w_STROBE_UMSB_0[11], w_STROBE_UMSB_0[10], w_STROBE_UMSB_0[9], w_STROBE_UMSB_0[8] } )
     );

UMSB_NB_INPUTS_4_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_8 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_umsb_2(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { w_umsb2_INPUTS[3], w_umsb2_INPUTS[2], w_umsb2_INPUTS[1], w_umsb2_INPUTS[0] } )
      , .OUTPUTS( { wire_INPUTS_0_11, wire_INPUTS_0_10, wire_INPUTS_0_9, wire_INPUTS_0_8 } )
      , .STROBE( { w_STROBE_UMSB_0[23], w_STROBE_UMSB_0[22], w_STROBE_UMSB_0[21], w_STROBE_UMSB_0[20], w_STROBE_UMSB_0[19], w_STROBE_UMSB_0[18], w_STROBE_UMSB_0[17], w_STROBE_UMSB_0[16] } )
     );

UMSB_NB_INPUTS_4_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_8 cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop_umsb_3(
        .DATA( { cluster_data1[7], cluster_data1[6], cluster_data1[5], cluster_data1[4], cluster_data1[3], cluster_data1[2], cluster_data1[1], cluster_data1[0] } )
      , .INPUTS( { w_umsb3_INPUTS[3], w_umsb3_INPUTS[2], w_umsb3_INPUTS[1], w_umsb3_INPUTS[0] } )
      , .OUTPUTS( { wire_INPUTS_0_15, wire_INPUTS_0_14, wire_INPUTS_0_13, wire_INPUTS_0_12 } )
      , .STROBE( { w_STROBE_UMSB_0[31], w_STROBE_UMSB_0[30], w_STROBE_UMSB_0[29], w_STROBE_UMSB_0[28], w_STROBE_UMSB_0[27], w_STROBE_UMSB_0[26], w_STROBE_UMSB_0[25], w_STROBE_UMSB_0[24] } )
     );

loader_type2_addressSize_9 loader_cluster_1_ins_cluster_l_1_TileBoundaryTop_TileBoundaryTop(
        .CLK( conf_ck1 )
      , .RESET( reset1 )
      , .SELECT_LEVEL( selector1 )
      , .ADDRESS( { address1[8], address1[7], address1[6], address1[5], address1[4], address1[3], address1[2], address1[1], address1[0] } )
      , .ADDRESS_LEVEL_D( { w_ADDRESS_LEVEL_D_0[5], w_ADDRESS_LEVEL_D_0[4], w_ADDRESS_LEVEL_D_0[3], w_ADDRESS_LEVEL_D_0[2], w_ADDRESS_LEVEL_D_0[1], w_ADDRESS_LEVEL_D_0[0] } )
      , .SELECT_LEVEL_D( { w_SELECT_LEVEL_D_0[3], w_SELECT_LEVEL_D_0[2], w_SELECT_LEVEL_D_0[1], w_SELECT_LEVEL_D_0[0] } )
      , .STROBE_DMSB( { w_STROBE_DMSB_0[63], w_STROBE_DMSB_0[62], w_STROBE_DMSB_0[61], w_STROBE_DMSB_0[60], w_STROBE_DMSB_0[59], w_STROBE_DMSB_0[58], w_STROBE_DMSB_0[57], w_STROBE_DMSB_0[56], w_STROBE_DMSB_0[55], w_STROBE_DMSB_0[54], w_STROBE_DMSB_0[53], w_STROBE_DMSB_0[52], w_STROBE_DMSB_0[51], w_STROBE_DMSB_0[50], w_STROBE_DMSB_0[49], w_STROBE_DMSB_0[48], w_STROBE_DMSB_0[47], w_STROBE_DMSB_0[46], w_STROBE_DMSB_0[45], w_STROBE_DMSB_0[44], w_STROBE_DMSB_0[43], w_STROBE_DMSB_0[42], w_STROBE_DMSB_0[41], w_STROBE_DMSB_0[40], w_STROBE_DMSB_0[39], w_STROBE_DMSB_0[38], w_STROBE_DMSB_0[37], w_STROBE_DMSB_0[36], w_STROBE_DMSB_0[35], w_STROBE_DMSB_0[34], w_STROBE_DMSB_0[33], w_STROBE_DMSB_0[32], w_STROBE_DMSB_0[31], w_STROBE_DMSB_0[30], w_STROBE_DMSB_0[29], w_STROBE_DMSB_0[28], w_STROBE_DMSB_0[27], w_STROBE_DMSB_0[26], w_STROBE_DMSB_0[25], w_STROBE_DMSB_0[24], w_STROBE_DMSB_0[23], w_STROBE_DMSB_0[22], w_STROBE_DMSB_0[21], w_STROBE_DMSB_0[20], w_STROBE_DMSB_0[19], w_STROBE_DMSB_0[18], w_STROBE_DMSB_0[17], w_STROBE_DMSB_0[16], w_STROBE_DMSB_0[15], w_STROBE_DMSB_0[14], w_STROBE_DMSB_0[13], w_STROBE_DMSB_0[12], w_STROBE_DMSB_0[11], w_STROBE_DMSB_0[10], w_STROBE_DMSB_0[9], w_STROBE_DMSB_0[8], w_STROBE_DMSB_0[7], w_STROBE_DMSB_0[6], w_STROBE_DMSB_0[5], w_STROBE_DMSB_0[4], w_STROBE_DMSB_0[3], w_STROBE_DMSB_0[2], w_STROBE_DMSB_0[1], w_STROBE_DMSB_0[0] } )
      , .STROBE_UMSB( { w_STROBE_UMSB_0[31], w_STROBE_UMSB_0[30], w_STROBE_UMSB_0[29], w_STROBE_UMSB_0[28], w_STROBE_UMSB_0[27], w_STROBE_UMSB_0[26], w_STROBE_UMSB_0[25], w_STROBE_UMSB_0[24], w_STROBE_UMSB_0[23], w_STROBE_UMSB_0[22], w_STROBE_UMSB_0[21], w_STROBE_UMSB_0[20], w_STROBE_UMSB_0[19], w_STROBE_UMSB_0[18], w_STROBE_UMSB_0[17], w_STROBE_UMSB_0[16], w_STROBE_UMSB_0[15], w_STROBE_UMSB_0[14], w_STROBE_UMSB_0[13], w_STROBE_UMSB_0[12], w_STROBE_UMSB_0[11], w_STROBE_UMSB_0[10], w_STROBE_UMSB_0[9], w_STROBE_UMSB_0[8], w_STROBE_UMSB_0[7], w_STROBE_UMSB_0[6], w_STROBE_UMSB_0[5], w_STROBE_UMSB_0[4], w_STROBE_UMSB_0[3], w_STROBE_UMSB_0[2], w_STROBE_UMSB_0[1], w_STROBE_UMSB_0[0] } )
     );


endmodule
