`timescale 1 ns/1 ps

module cluster_0(
     func_ck0
   , conf_ck0
   , selector0
   , reset0
   , input_tree0
   , output_tree0
   , cluster_inputs0
   , cluster_outputs0
   , cluster_data0
   , address0
  );


input   func_ck0;
wire func_ck0;
input   conf_ck0;
wire conf_ck0;
input   selector0;
wire selector0;
input   reset0;
wire reset0;
input   [15:0] input_tree0;
wire [15:0] input_tree0;
output  [3:0] output_tree0;
wire [3:0] output_tree0;
input   [15:0] cluster_inputs0;
wire [15:0] cluster_inputs0;
output  [3:0] cluster_outputs0;
wire [3:0] cluster_outputs0;
input   [7:0] cluster_data0;
wire [7:0] cluster_data0;
input   [5:0] address0;
wire [5:0] address0;

wire wire_OUTPUTS_4_0;
wire wire_OUTPUTS_4_1;
wire wire_OUTPUTS_4_2;
wire wire_OUTPUTS_4_3;
wire wire_STROBE_0_0;
wire wire_STROBE_10_0;
wire wire_STROBE_11_0;
wire wire_STROBE_12_0;
wire wire_STROBE_13_0;
wire wire_STROBE_14_0;
wire wire_STROBE_15_0;
wire wire_STROBE_16_0;
wire wire_STROBE_17_0;
wire wire_STROBE_18_0;
wire wire_STROBE_19_0;
wire wire_STROBE_1_0;
wire wire_STROBE_2_0;
wire wire_STROBE_3_0;
wire wire_STROBE_4_0;
wire wire_STROBE_5_0;
wire wire_STROBE_6_0;
wire wire_STROBE_7_0;
wire wire_STROBE_8_0;
wire wire_STROBE_9_0;
wire [67:0] w_STROBE_BLE_0;
wire [7:0] w_STROBE_DMSBOUT_0;
wire [59:0] w_STROBE_DMSB_0;
wire [3:0] w_dmsb0_OUTPUTS;
wire [3:0] w_dmsb1_OUTPUTS;
wire [3:0] w_dmsb2_OUTPUTS;
wire [3:0] w_dmsb3_OUTPUTS;
wire [3:0] w_umsb0_INPUTS;

BLE_NB_INPUTS_4_DATA_SIZE_8 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_ble_0(
        .CLK( func_ck0 )
      , .OUTPUT( w_umsb0_INPUTS[0] )
      , .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { w_dmsb3_OUTPUTS[0], w_dmsb2_OUTPUTS[0], w_dmsb1_OUTPUTS[0], w_dmsb0_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_BLE_0[16], w_STROBE_BLE_0[15], w_STROBE_BLE_0[14], w_STROBE_BLE_0[13], w_STROBE_BLE_0[12], w_STROBE_BLE_0[11], w_STROBE_BLE_0[10], w_STROBE_BLE_0[9], w_STROBE_BLE_0[8], w_STROBE_BLE_0[7], w_STROBE_BLE_0[6], w_STROBE_BLE_0[5], w_STROBE_BLE_0[4], w_STROBE_BLE_0[3], w_STROBE_BLE_0[2], w_STROBE_BLE_0[1], w_STROBE_BLE_0[0] } )
     );

BLE_NB_INPUTS_4_DATA_SIZE_8 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_ble_1(
        .CLK( func_ck0 )
      , .OUTPUT( w_umsb0_INPUTS[1] )
      , .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { w_dmsb3_OUTPUTS[1], w_dmsb2_OUTPUTS[1], w_dmsb1_OUTPUTS[1], w_dmsb0_OUTPUTS[1] } )
      , .STROBE( { w_STROBE_BLE_0[33], w_STROBE_BLE_0[32], w_STROBE_BLE_0[31], w_STROBE_BLE_0[30], w_STROBE_BLE_0[29], w_STROBE_BLE_0[28], w_STROBE_BLE_0[27], w_STROBE_BLE_0[26], w_STROBE_BLE_0[25], w_STROBE_BLE_0[24], w_STROBE_BLE_0[23], w_STROBE_BLE_0[22], w_STROBE_BLE_0[21], w_STROBE_BLE_0[20], w_STROBE_BLE_0[19], w_STROBE_BLE_0[18], w_STROBE_BLE_0[17] } )
     );

BLE_NB_INPUTS_4_DATA_SIZE_8 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_ble_2(
        .CLK( func_ck0 )
      , .OUTPUT( w_umsb0_INPUTS[2] )
      , .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { w_dmsb3_OUTPUTS[2], w_dmsb2_OUTPUTS[2], w_dmsb1_OUTPUTS[2], w_dmsb0_OUTPUTS[2] } )
      , .STROBE( { w_STROBE_BLE_0[50], w_STROBE_BLE_0[49], w_STROBE_BLE_0[48], w_STROBE_BLE_0[47], w_STROBE_BLE_0[46], w_STROBE_BLE_0[45], w_STROBE_BLE_0[44], w_STROBE_BLE_0[43], w_STROBE_BLE_0[42], w_STROBE_BLE_0[41], w_STROBE_BLE_0[40], w_STROBE_BLE_0[39], w_STROBE_BLE_0[38], w_STROBE_BLE_0[37], w_STROBE_BLE_0[36], w_STROBE_BLE_0[35], w_STROBE_BLE_0[34] } )
     );

BLE_NB_INPUTS_4_DATA_SIZE_8 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_ble_3(
        .CLK( func_ck0 )
      , .OUTPUT( w_umsb0_INPUTS[3] )
      , .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { w_dmsb3_OUTPUTS[3], w_dmsb2_OUTPUTS[3], w_dmsb1_OUTPUTS[3], w_dmsb0_OUTPUTS[3] } )
      , .STROBE( { w_STROBE_BLE_0[67], w_STROBE_BLE_0[66], w_STROBE_BLE_0[65], w_STROBE_BLE_0[64], w_STROBE_BLE_0[63], w_STROBE_BLE_0[62], w_STROBE_BLE_0[61], w_STROBE_BLE_0[60], w_STROBE_BLE_0[59], w_STROBE_BLE_0[58], w_STROBE_BLE_0[57], w_STROBE_BLE_0[56], w_STROBE_BLE_0[55], w_STROBE_BLE_0[54], w_STROBE_BLE_0[53], w_STROBE_BLE_0[52], w_STROBE_BLE_0[51] } )
     );

DMSB_NB_INPUTS_5_DATA_SIZE_8_NB_OUTPUTS_5_STROBE_SIZE_15 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_dmsb_0(
        .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { cluster_outputs0[0], cluster_inputs0[3], cluster_inputs0[2], cluster_inputs0[1], cluster_inputs0[0] } )
      , .OUTPUTS( { wire_OUTPUTS_4_0, w_dmsb0_OUTPUTS[3], w_dmsb0_OUTPUTS[2], w_dmsb0_OUTPUTS[1], w_dmsb0_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[14], w_STROBE_DMSB_0[13], w_STROBE_DMSB_0[12], w_STROBE_DMSB_0[11], w_STROBE_DMSB_0[10], w_STROBE_DMSB_0[9], w_STROBE_DMSB_0[8], w_STROBE_DMSB_0[7], w_STROBE_DMSB_0[6], w_STROBE_DMSB_0[5], w_STROBE_DMSB_0[4], w_STROBE_DMSB_0[3], w_STROBE_DMSB_0[2], w_STROBE_DMSB_0[1], w_STROBE_DMSB_0[0] } )
     );

DMSB_NB_INPUTS_5_DATA_SIZE_8_NB_OUTPUTS_5_STROBE_SIZE_15 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_dmsb_1(
        .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { cluster_outputs0[1], cluster_inputs0[7], cluster_inputs0[6], cluster_inputs0[5], cluster_inputs0[4] } )
      , .OUTPUTS( { wire_OUTPUTS_4_1, w_dmsb1_OUTPUTS[3], w_dmsb1_OUTPUTS[2], w_dmsb1_OUTPUTS[1], w_dmsb1_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[29], w_STROBE_DMSB_0[28], w_STROBE_DMSB_0[27], w_STROBE_DMSB_0[26], w_STROBE_DMSB_0[25], w_STROBE_DMSB_0[24], w_STROBE_DMSB_0[23], w_STROBE_DMSB_0[22], w_STROBE_DMSB_0[21], w_STROBE_DMSB_0[20], w_STROBE_DMSB_0[19], w_STROBE_DMSB_0[18], w_STROBE_DMSB_0[17], w_STROBE_DMSB_0[16], w_STROBE_DMSB_0[15] } )
     );

DMSB_NB_INPUTS_5_DATA_SIZE_8_NB_OUTPUTS_5_STROBE_SIZE_15 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_dmsb_2(
        .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { cluster_outputs0[2], cluster_inputs0[11], cluster_inputs0[10], cluster_inputs0[9], cluster_inputs0[8] } )
      , .OUTPUTS( { wire_OUTPUTS_4_2, w_dmsb2_OUTPUTS[3], w_dmsb2_OUTPUTS[2], w_dmsb2_OUTPUTS[1], w_dmsb2_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[44], w_STROBE_DMSB_0[43], w_STROBE_DMSB_0[42], w_STROBE_DMSB_0[41], w_STROBE_DMSB_0[40], w_STROBE_DMSB_0[39], w_STROBE_DMSB_0[38], w_STROBE_DMSB_0[37], w_STROBE_DMSB_0[36], w_STROBE_DMSB_0[35], w_STROBE_DMSB_0[34], w_STROBE_DMSB_0[33], w_STROBE_DMSB_0[32], w_STROBE_DMSB_0[31], w_STROBE_DMSB_0[30] } )
     );

DMSB_NB_INPUTS_5_DATA_SIZE_8_NB_OUTPUTS_5_STROBE_SIZE_15 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_dmsb_3(
        .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { cluster_outputs0[3], cluster_inputs0[15], cluster_inputs0[14], cluster_inputs0[13], cluster_inputs0[12] } )
      , .OUTPUTS( { wire_OUTPUTS_4_3, w_dmsb3_OUTPUTS[3], w_dmsb3_OUTPUTS[2], w_dmsb3_OUTPUTS[1], w_dmsb3_OUTPUTS[0] } )
      , .STROBE( { w_STROBE_DMSB_0[59], w_STROBE_DMSB_0[58], w_STROBE_DMSB_0[57], w_STROBE_DMSB_0[56], w_STROBE_DMSB_0[55], w_STROBE_DMSB_0[54], w_STROBE_DMSB_0[53], w_STROBE_DMSB_0[52], w_STROBE_DMSB_0[51], w_STROBE_DMSB_0[50], w_STROBE_DMSB_0[49], w_STROBE_DMSB_0[48], w_STROBE_DMSB_0[47], w_STROBE_DMSB_0[46], w_STROBE_DMSB_0[45] } )
     );

DMSB_NB_INPUTS_4_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_8 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_dmsbout(
        .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { wire_OUTPUTS_4_3, wire_OUTPUTS_4_2, wire_OUTPUTS_4_1, wire_OUTPUTS_4_0 } )
      , .OUTPUTS( { output_tree0[3], output_tree0[2], output_tree0[1], output_tree0[0] } )
      , .STROBE( { w_STROBE_DMSBOUT_0[7], w_STROBE_DMSBOUT_0[6], w_STROBE_DMSBOUT_0[5], w_STROBE_DMSBOUT_0[4], w_STROBE_DMSBOUT_0[3], w_STROBE_DMSBOUT_0[2], w_STROBE_DMSBOUT_0[1], w_STROBE_DMSBOUT_0[0] } )
     );

UMSB_NB_INPUTS_20_DATA_SIZE_8_NB_OUTPUTS_4_STROBE_SIZE_20 cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop_umsb_0(
        .DATA( { cluster_data0[7], cluster_data0[6], cluster_data0[5], cluster_data0[4], cluster_data0[3], cluster_data0[2], cluster_data0[1], cluster_data0[0] } )
      , .INPUTS( { input_tree0[15], input_tree0[14], input_tree0[13], input_tree0[12], input_tree0[11], input_tree0[10], input_tree0[9], input_tree0[8], input_tree0[7], input_tree0[6], input_tree0[5], input_tree0[4], input_tree0[3], input_tree0[2], input_tree0[1], input_tree0[0], w_umsb0_INPUTS[3], w_umsb0_INPUTS[2], w_umsb0_INPUTS[1], w_umsb0_INPUTS[0] } )
      , .OUTPUTS( { cluster_outputs0[3], cluster_outputs0[2], cluster_outputs0[1], cluster_outputs0[0] } )
      , .STROBE( { wire_STROBE_19_0, wire_STROBE_18_0, wire_STROBE_17_0, wire_STROBE_16_0, wire_STROBE_15_0, wire_STROBE_14_0, wire_STROBE_13_0, wire_STROBE_12_0, wire_STROBE_11_0, wire_STROBE_10_0, wire_STROBE_9_0, wire_STROBE_8_0, wire_STROBE_7_0, wire_STROBE_6_0, wire_STROBE_5_0, wire_STROBE_4_0, wire_STROBE_3_0, wire_STROBE_2_0, wire_STROBE_1_0, wire_STROBE_0_0 } )
     );

loader_0_addressSize_6 loader_cluster_0_instance_cluster0_TileBoundaryTop_TileBoundaryTop(
        .CLK( conf_ck0 )
      , .RESET( reset0 )
      , .SELECT_LEVEL( selector0 )
      , .ADDRESS( { address0[5], address0[4], address0[3], address0[2], address0[1], address0[0] } )
      , .STROBE_BLE( { w_STROBE_BLE_0[67], w_STROBE_BLE_0[66], w_STROBE_BLE_0[65], w_STROBE_BLE_0[64], w_STROBE_BLE_0[63], w_STROBE_BLE_0[62], w_STROBE_BLE_0[61], w_STROBE_BLE_0[60], w_STROBE_BLE_0[59], w_STROBE_BLE_0[58], w_STROBE_BLE_0[57], w_STROBE_BLE_0[56], w_STROBE_BLE_0[55], w_STROBE_BLE_0[54], w_STROBE_BLE_0[53], w_STROBE_BLE_0[52], w_STROBE_BLE_0[51], w_STROBE_BLE_0[50], w_STROBE_BLE_0[49], w_STROBE_BLE_0[48], w_STROBE_BLE_0[47], w_STROBE_BLE_0[46], w_STROBE_BLE_0[45], w_STROBE_BLE_0[44], w_STROBE_BLE_0[43], w_STROBE_BLE_0[42], w_STROBE_BLE_0[41], w_STROBE_BLE_0[40], w_STROBE_BLE_0[39], w_STROBE_BLE_0[38], w_STROBE_BLE_0[37], w_STROBE_BLE_0[36], w_STROBE_BLE_0[35], w_STROBE_BLE_0[34], w_STROBE_BLE_0[33], w_STROBE_BLE_0[32], w_STROBE_BLE_0[31], w_STROBE_BLE_0[30], w_STROBE_BLE_0[29], w_STROBE_BLE_0[28], w_STROBE_BLE_0[27], w_STROBE_BLE_0[26], w_STROBE_BLE_0[25], w_STROBE_BLE_0[24], w_STROBE_BLE_0[23], w_STROBE_BLE_0[22], w_STROBE_BLE_0[21], w_STROBE_BLE_0[20], w_STROBE_BLE_0[19], w_STROBE_BLE_0[18], w_STROBE_BLE_0[17], w_STROBE_BLE_0[16], w_STROBE_BLE_0[15], w_STROBE_BLE_0[14], w_STROBE_BLE_0[13], w_STROBE_BLE_0[12], w_STROBE_BLE_0[11], w_STROBE_BLE_0[10], w_STROBE_BLE_0[9], w_STROBE_BLE_0[8], w_STROBE_BLE_0[7], w_STROBE_BLE_0[6], w_STROBE_BLE_0[5], w_STROBE_BLE_0[4], w_STROBE_BLE_0[3], w_STROBE_BLE_0[2], w_STROBE_BLE_0[1], w_STROBE_BLE_0[0] } )
      , .STROBE_DMSB( { w_STROBE_DMSB_0[59], w_STROBE_DMSB_0[58], w_STROBE_DMSB_0[57], w_STROBE_DMSB_0[56], w_STROBE_DMSB_0[55], w_STROBE_DMSB_0[54], w_STROBE_DMSB_0[53], w_STROBE_DMSB_0[52], w_STROBE_DMSB_0[51], w_STROBE_DMSB_0[50], w_STROBE_DMSB_0[49], w_STROBE_DMSB_0[48], w_STROBE_DMSB_0[47], w_STROBE_DMSB_0[46], w_STROBE_DMSB_0[45], w_STROBE_DMSB_0[44], w_STROBE_DMSB_0[43], w_STROBE_DMSB_0[42], w_STROBE_DMSB_0[41], w_STROBE_DMSB_0[40], w_STROBE_DMSB_0[39], w_STROBE_DMSB_0[38], w_STROBE_DMSB_0[37], w_STROBE_DMSB_0[36], w_STROBE_DMSB_0[35], w_STROBE_DMSB_0[34], w_STROBE_DMSB_0[33], w_STROBE_DMSB_0[32], w_STROBE_DMSB_0[31], w_STROBE_DMSB_0[30], w_STROBE_DMSB_0[29], w_STROBE_DMSB_0[28], w_STROBE_DMSB_0[27], w_STROBE_DMSB_0[26], w_STROBE_DMSB_0[25], w_STROBE_DMSB_0[24], w_STROBE_DMSB_0[23], w_STROBE_DMSB_0[22], w_STROBE_DMSB_0[21], w_STROBE_DMSB_0[20], w_STROBE_DMSB_0[19], w_STROBE_DMSB_0[18], w_STROBE_DMSB_0[17], w_STROBE_DMSB_0[16], w_STROBE_DMSB_0[15], w_STROBE_DMSB_0[14], w_STROBE_DMSB_0[13], w_STROBE_DMSB_0[12], w_STROBE_DMSB_0[11], w_STROBE_DMSB_0[10], w_STROBE_DMSB_0[9], w_STROBE_DMSB_0[8], w_STROBE_DMSB_0[7], w_STROBE_DMSB_0[6], w_STROBE_DMSB_0[5], w_STROBE_DMSB_0[4], w_STROBE_DMSB_0[3], w_STROBE_DMSB_0[2], w_STROBE_DMSB_0[1], w_STROBE_DMSB_0[0] } )
      , .STROBE_DMSBOUT( { w_STROBE_DMSBOUT_0[7], w_STROBE_DMSBOUT_0[6], w_STROBE_DMSBOUT_0[5], w_STROBE_DMSBOUT_0[4], w_STROBE_DMSBOUT_0[3], w_STROBE_DMSBOUT_0[2], w_STROBE_DMSBOUT_0[1], w_STROBE_DMSBOUT_0[0] } )
      , .STROBE_UMSB( { wire_STROBE_19_0, wire_STROBE_18_0, wire_STROBE_17_0, wire_STROBE_16_0, wire_STROBE_15_0, wire_STROBE_14_0, wire_STROBE_13_0, wire_STROBE_12_0, wire_STROBE_11_0, wire_STROBE_10_0, wire_STROBE_9_0, wire_STROBE_8_0, wire_STROBE_7_0, wire_STROBE_6_0, wire_STROBE_5_0, wire_STROBE_4_0, wire_STROBE_3_0, wire_STROBE_2_0, wire_STROBE_1_0, wire_STROBE_0_0 } )
     );


endmodule
